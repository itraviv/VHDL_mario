--------------------------------------
-- SinTable.vhd
-- Written by Saar Eliad and Itamar Raviv.
-- All rights reserved, Copyright 2017
--------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity BombSoundTable is
port(
  CLK     : in std_logic;
  RESET_N : in std_logic;
  ENA     : in std_logic;
  ADDR    : in std_logic_vector(11 downto 0);
  Q       : out std_logic_vector(7 downto 0)
);
end BombSoundTable;

architecture arch of BombSoundTable is

type table_type is array(0 to 4095) of std_logic_vector(7 downto 0);
signal sqr_table : table_type;

begin

  BombSoundTable_proc: process(RESET_N, CLK)
    constant sqr_table : table_type := (
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FE",
X"F0",
X"FB",
X"04",
X"16",
X"00",
X"F9",
X"07",
X"FF",
X"07",
X"07",
X"0C",
X"0C",
X"16",
X"0B",
X"00",
X"09",
X"09",
X"F6",
X"FC",
X"E9",
X"E3",
X"F0",
X"F8",
X"FF",
X"E4",
X"00",
X"03",
X"FC",
X"06",
X"F5",
X"04",
X"0F",
X"FE",
X"00",
X"09",
X"F5",
X"00",
X"07",
X"06",
X"00",
X"02",
X"22",
X"26",
X"D6",
X"E7",
X"0A",
X"35",
X"0D",
X"F9",
X"D6",
X"E1",
X"11",
X"C7",
X"F4",
X"D6",
X"00",
X"01",
X"EA",
X"DF",
X"00",
X"EE",
X"FD",
X"FA",
X"09",
X"0E",
X"03",
X"0E",
X"EF",
X"1E",
X"00",
X"02",
X"03",
X"13",
X"0A",
X"FF",
X"FE",
X"1A",
X"00",
X"0E",
X"1E",
X"0D",
X"1F",
X"0E",
X"15",
X"10",
X"FC",
X"05",
X"FB",
X"09",
X"01",
X"F6",
X"E7",
X"06",
X"F2",
X"FB",
X"03",
X"F9",
X"0C",
X"DC",
X"FF",
X"00",
X"E4",
X"DB",
X"F5",
X"DE",
X"FC",
X"E4",
X"FD",
X"EB",
X"EA",
X"E4",
X"FF",
X"FE",
X"FA",
X"16",
X"0C",
X"24",
X"00",
X"1E",
X"00",
X"14",
X"0A",
X"19",
X"18",
X"0A",
X"02",
X"F4",
X"0C",
X"03",
X"FF",
X"0B",
X"FA",
X"FF",
X"09",
X"FA",
X"FC",
X"F2",
X"F3",
X"EC",
X"FE",
X"E8",
X"FD",
X"EA",
X"00",
X"E1",
X"F0",
X"08",
X"40",
X"F9",
X"CA",
X"0A",
X"14",
X"19",
X"EB",
X"1C",
X"00",
X"15",
X"3A",
X"1A",
X"FF",
X"D2",
X"38",
X"15",
X"F8",
X"21",
X"EE",
X"43",
X"1C",
X"FA",
X"32",
X"06",
X"E1",
X"F2",
X"1D",
X"E6",
X"16",
X"EB",
X"C2",
X"0F",
X"C2",
X"F8",
X"D6",
X"CD",
X"E6",
X"D6",
X"CF",
X"C5",
X"0E",
X"B3",
X"06",
X"E4",
X"E1",
X"25",
X"BE",
X"10",
X"0E",
X"E9",
X"31",
X"07",
X"EB",
X"25",
X"F5",
X"19",
X"20",
X"12",
X"2A",
X"FF",
X"FE",
X"29",
X"28",
X"26",
X"20",
X"15",
X"21",
X"08",
X"1C",
X"11",
X"03",
X"20",
X"03",
X"05",
X"00",
X"06",
X"01",
X"06",
X"00",
X"00",
X"F2",
X"E9",
X"E8",
X"06",
X"BB",
X"DF",
X"DF",
X"AE",
X"BA",
X"CE",
X"D8",
X"F4",
X"F4",
X"10",
X"1C",
X"F9",
X"ED",
X"BB",
X"CE",
X"EC",
X"06",
X"04",
X"1F",
X"0B",
X"2E",
X"1E",
X"14",
X"FF",
X"00",
X"1C",
X"2A",
X"26",
X"2B",
X"2B",
X"F1",
X"03",
X"13",
X"18",
X"1A",
X"32",
X"3C",
X"F8",
X"D6",
X"F7",
X"25",
X"FA",
X"DA",
X"F6",
X"0D",
X"F3",
X"D7",
X"EA",
X"0B",
X"FA",
X"14",
X"19",
X"15",
X"31",
X"DC",
X"F6",
X"DE",
X"03",
X"E1",
X"E3",
X"E2",
X"E2",
X"E9",
X"D7",
X"F1",
X"EC",
X"0A",
X"DE",
X"06",
X"13",
X"E4",
X"EC",
X"EA",
X"F7",
X"E5",
X"DD",
X"C8",
X"06",
X"0B",
X"11",
X"07",
X"10",
X"09",
X"35",
X"28",
X"37",
X"35",
X"2C",
X"1D",
X"43",
X"29",
X"1F",
X"F4",
X"1E",
X"04",
X"13",
X"FE",
X"DB",
X"12",
X"E6",
X"EB",
X"01",
X"22",
X"D5",
X"03",
X"FC",
X"24",
X"E4",
X"09",
X"F1",
X"D9",
X"ED",
X"F6",
X"C3",
X"F5",
X"D0",
X"C8",
X"0E",
X"CD",
X"EE",
X"0A",
X"DB",
X"DE",
X"23",
X"FE",
X"05",
X"06",
X"F0",
X"00",
X"00",
X"FD",
X"C9",
X"F8",
X"C7",
X"0B",
X"2D",
X"EC",
X"0E",
X"51",
X"11",
X"06",
X"64",
X"52",
X"0B",
X"4F",
X"04",
X"36",
X"1B",
X"00",
X"0E",
X"01",
X"0C",
X"EA",
X"05",
X"05",
X"F2",
X"00",
X"FA",
X"FC",
X"E6",
X"F2",
X"E6",
X"D3",
X"E9",
X"CD",
X"03",
X"06",
X"E6",
X"E0",
X"E1",
X"DC",
X"DF",
X"EC",
X"E8",
X"ED",
X"FD",
X"E4",
X"D9",
X"FB",
X"0E",
X"E2",
X"F2",
X"3E",
X"F5",
X"30",
X"1E",
X"10",
X"29",
X"25",
X"43",
X"24",
X"1E",
X"3E",
X"03",
X"FE",
X"15",
X"D0",
X"FF",
X"E8",
X"F7",
X"E9",
X"E6",
X"0A",
X"03",
X"D9",
X"F5",
X"03",
X"E5",
X"13",
X"0B",
X"EC",
X"08",
X"1F",
X"33",
X"FD",
X"06",
X"11",
X"E9",
X"DE",
X"FC",
X"C3",
X"E8",
X"F5",
X"07",
X"00",
X"11",
X"00",
X"11",
X"F6",
X"1C",
X"0A",
X"FB",
X"FB",
X"E5",
X"E7",
X"0B",
X"FF",
X"1D",
X"12",
X"19",
X"09",
X"EF",
X"F2",
X"E4",
X"DF",
X"D9",
X"E2",
X"DF",
X"C2",
X"04",
X"1A",
X"E2",
X"02",
X"1A",
X"40",
X"28",
X"FB",
X"31",
X"38",
X"0E",
X"28",
X"FA",
X"05",
X"33",
X"12",
X"00",
X"FB",
X"F5",
X"C2",
X"06",
X"EA",
X"CC",
X"03",
X"07",
X"00",
X"19",
X"08",
X"F4",
X"FC",
X"02",
X"DD",
X"F1",
X"F5",
X"E5",
X"FD",
X"03",
X"FA",
X"09",
X"1B",
X"02",
X"11",
X"C6",
X"00",
X"E7",
X"17",
X"BD",
X"E3",
X"06",
X"E0",
X"14",
X"09",
X"D0",
X"12",
X"E5",
X"DB",
X"0D",
X"F7",
X"F2",
X"4B",
X"05",
X"24",
X"0D",
X"1E",
X"27",
X"29",
X"0B",
X"1E",
X"14",
X"1C",
X"27",
X"08",
X"14",
X"FE",
X"15",
X"01",
X"04",
X"F2",
X"00",
X"E9",
X"F9",
X"DD",
X"F2",
X"E5",
X"DE",
X"EC",
X"EE",
X"EC",
X"E7",
X"E1",
X"F2",
X"F1",
X"F1",
X"EB",
X"0D",
X"EC",
X"E7",
X"00",
X"F6",
X"0A",
X"00",
X"19",
X"0D",
X"1F",
X"21",
X"0D",
X"FF",
X"0A",
X"0D",
X"00",
X"04",
X"FA",
X"05",
X"05",
X"F3",
X"FB",
X"0E",
X"16",
X"FB",
X"FA",
X"15",
X"10",
X"F9",
X"F2",
X"11",
X"03",
X"18",
X"EF",
X"08",
X"16",
X"E9",
X"0B",
X"00",
X"03",
X"29",
X"09",
X"FC",
X"0A",
X"F7",
X"01",
X"F5",
X"E5",
X"ED",
X"E4",
X"EA",
X"E2",
X"FB",
X"E7",
X"EA",
X"F8",
X"EE",
X"04",
X"F6",
X"F9",
X"0F",
X"F8",
X"00",
X"FA",
X"FE",
X"03",
X"EE",
X"FC",
X"00",
X"05",
X"09",
X"10",
X"0D",
X"12",
X"12",
X"FD",
X"14",
X"FE",
X"29",
X"04",
X"03",
X"14",
X"01",
X"1F",
X"11",
X"15",
X"EC",
X"DF",
X"11",
X"ED",
X"F0",
X"04",
X"FB",
X"F4",
X"F4",
X"F3",
X"F8",
X"EC",
X"11",
X"DC",
X"D3",
X"F0",
X"F6",
X"F6",
X"F0",
X"02",
X"FD",
X"FC",
X"F2",
X"02",
X"02",
X"0E",
X"1E",
X"EE",
X"EE",
X"0D",
X"01",
X"05",
X"03",
X"21",
X"07",
X"F1",
X"01",
X"01",
X"29",
X"03",
X"04",
X"04",
X"EF",
X"00",
X"FF",
X"F8",
X"11",
X"14",
X"02",
X"21",
X"0F",
X"FD",
X"2B",
X"26",
X"F2",
X"E4",
X"F3",
X"0F",
X"F8",
X"00",
X"0E",
X"08",
X"FB",
X"F8",
X"E2",
X"EB",
X"E2",
X"E4",
X"D5",
X"E3",
X"DE",
X"EA",
X"F9",
X"EB",
X"F7",
X"F5",
X"FE",
X"F3",
X"F6",
X"F7",
X"16",
X"1F",
X"09",
X"09",
X"0D",
X"29",
X"21",
X"10",
X"20",
X"15",
X"18",
X"FE",
X"16",
X"00",
X"ED",
X"0E",
X"FB",
X"F7",
X"00",
X"05",
X"DE",
X"FF",
X"00",
X"23",
X"F9",
X"00",
X"06",
X"11",
X"FA",
X"04",
X"05",
X"03",
X"00",
X"02",
X"F1",
X"F3",
X"F7",
X"F0",
X"E4",
X"E3",
X"DB",
X"D4",
X"D4",
X"F2",
X"E1",
X"D9",
X"F3",
X"F2",
X"01",
X"0E",
X"09",
X"2C",
X"1A",
X"0C",
X"3A",
X"08",
X"1C",
X"17",
X"14",
X"12",
X"08",
X"04",
X"06",
X"05",
X"07",
X"0E",
X"0D",
X"19",
X"29",
X"10",
X"1F",
X"09",
X"17",
X"CF",
X"D2",
X"F4",
X"00",
X"FD",
X"FA",
X"F2",
X"ED",
X"E5",
X"D3",
X"D5",
X"D1",
X"D6",
X"D6",
X"D6",
X"E9",
X"07",
X"05",
X"00",
X"0F",
X"11",
X"0B",
X"0F",
X"0B",
X"07",
X"0A",
X"0C",
X"0A",
X"13",
X"11",
X"14",
X"12",
X"10",
X"0E",
X"0F",
X"0C",
X"0C",
X"08",
X"0A",
X"0F",
X"E6",
X"F0",
X"FA",
X"01",
X"07",
X"05",
X"00",
X"F8",
X"F6",
X"F3",
X"F1",
X"EF",
X"F3",
X"03",
X"08",
X"FF",
X"FC",
X"F9",
X"FD",
X"FB",
X"01",
X"0B",
X"0D",
X"08",
X"03",
X"FC",
X"F0",
X"E9",
X"E5",
X"DF",
X"DB",
X"DA",
X"DD",
X"DD",
X"E4",
X"EF",
X"F7",
X"02",
X"16",
X"1E",
X"2B",
X"35",
X"40",
X"45",
X"4B",
X"4C",
X"47",
X"3E",
X"34",
X"26",
X"17",
X"07",
X"F9",
X"E9",
X"DC",
X"CF",
X"C3",
X"B9",
X"B6",
X"B0",
X"B1",
X"B2",
X"BD",
X"C0",
X"BE",
X"D6",
X"DF",
X"FE",
X"08",
X"FE",
X"0C",
X"18",
X"21",
X"27",
X"1E",
X"2A",
X"2A",
X"27",
X"43",
X"43",
X"43",
X"39",
X"32",
X"24",
X"17",
X"0B",
X"08",
X"01",
X"F9",
X"F3",
X"F8",
X"FD",
X"EE",
X"E2",
X"E6",
X"EA",
X"E1",
X"F2",
X"FA",
X"E3",
X"DC",
X"D6",
X"D0",
X"D3",
X"D2",
X"DA",
X"DF",
X"E8",
X"F3",
X"FF",
X"03",
X"0E",
X"13",
X"1A",
X"20",
X"27",
X"27",
X"28",
X"21",
X"1B",
X"17",
X"12",
X"0D",
X"0D",
X"0A",
X"0E",
X"0B",
X"10",
X"0D",
X"0E",
X"06",
X"0C",
X"FF",
X"06",
X"FB",
X"EE",
X"F1",
X"DA",
X"D8",
X"E6",
X"E2",
X"DD",
X"DD",
X"E2",
X"E3",
X"DB",
X"D6",
X"F4",
X"10",
X"10",
X"19",
X"0A",
X"0F",
X"ED",
X"13",
X"00",
X"F0",
X"00",
X"03",
X"0F",
X"16",
X"17",
X"3A",
X"0C",
X"1A",
X"18",
X"11",
X"29",
X"08",
X"FD",
X"EA",
X"E9",
X"D0",
X"DA",
X"D8",
X"E5",
X"00",
X"0F",
X"13",
X"1A",
X"12",
X"0D",
X"FF",
X"F7",
X"F3",
X"F1",
X"F5",
X"FD",
X"FC",
X"08",
X"0D",
X"1F",
X"1B",
X"3A",
X"31",
X"14",
X"1F",
X"1D",
X"10",
X"01",
X"FB",
X"E9",
X"E2",
X"CF",
X"D9",
X"C4",
X"BF",
X"C6",
X"BE",
X"C3",
X"E0",
X"D5",
X"C6",
X"C7",
X"CE",
X"D8",
X"EE",
X"06",
X"1B",
X"2A",
X"3C",
X"40",
X"48",
X"4F",
X"3F",
X"30",
X"2A",
X"01",
X"10",
X"28",
X"FB",
X"0D",
X"35",
X"08",
X"15",
X"FE",
X"0C",
X"26",
X"F4",
X"32",
X"1E",
X"2C",
X"1E",
X"DF",
X"00",
X"02",
X"1F",
X"F5",
X"C4",
X"D1",
X"B8",
X"B9",
X"B2",
X"B4",
X"AF",
X"C4",
X"C7",
X"C7",
X"D3",
X"DD",
X"DA",
X"EE",
X"F8",
X"FF",
X"FD",
X"12",
X"26",
X"38",
X"20",
X"30",
X"3D",
X"22",
X"2C",
X"2F",
X"2A",
X"2A",
X"28",
X"1C",
X"15",
X"1D",
X"2B",
X"19",
X"18",
X"11",
X"FC",
X"FD",
X"FD",
X"F3",
X"E7",
X"DF",
X"DA",
X"DC",
X"DA",
X"D8",
X"E5",
X"F4",
X"EF",
X"E5",
X"F2",
X"F2",
X"00",
X"EC",
X"11",
X"DC",
X"E4",
X"FB",
X"00",
X"09",
X"05",
X"0D",
X"07",
X"0B",
X"12",
X"09",
X"12",
X"08",
X"00",
X"0A",
X"21",
X"25",
X"04",
X"00",
X"00",
X"08",
X"0A",
X"0D",
X"F8",
X"F0",
X"E2",
X"DC",
X"DF",
X"E3",
X"DD",
X"F6",
X"0B",
X"0E",
X"0F",
X"15",
X"1D",
X"20",
X"24",
X"1D",
X"17",
X"23",
X"0D",
X"0B",
X"DF",
X"E2",
X"E9",
X"D9",
X"EA",
X"DD",
X"CF",
X"CD",
X"BB",
X"D5",
X"EB",
X"DD",
X"FB",
X"23",
X"2D",
X"2A",
X"44",
X"2E",
X"36",
X"2F",
X"1D",
X"10",
X"1A",
X"0E",
X"F3",
X"10",
X"16",
X"14",
X"00",
X"01",
X"00",
X"EE",
X"F4",
X"F1",
X"EE",
X"EE",
X"EB",
X"EA",
X"E6",
X"E4",
X"E0",
X"DF",
X"E1",
X"DE",
X"E1",
X"E2",
X"DB",
X"E3",
X"EB",
X"F2",
X"F6",
X"F6",
X"FD",
X"03",
X"07",
X"14",
X"19",
X"24",
X"23",
X"34",
X"2C",
X"25",
X"1B",
X"1F",
X"16",
X"2A",
X"FC",
X"1E",
X"28",
X"04",
X"24",
X"18",
X"1B",
X"0A",
X"00",
X"F5",
X"EC",
X"DA",
X"C0",
X"C6",
X"EE",
X"DA",
X"BC",
X"C5",
X"B1",
X"B6",
X"CE",
X"E1",
X"FA",
X"05",
X"11",
X"14",
X"0F",
X"0C",
X"0B",
X"1B",
X"0E",
X"04",
X"14",
X"0F",
X"08",
X"00",
X"0A",
X"14",
X"1A",
X"2D",
X"2F",
X"33",
X"2B",
X"2C",
X"30",
X"2A",
X"29",
X"1C",
X"20",
X"04",
X"03",
X"00",
X"EE",
X"E3",
X"D0",
X"D0",
X"D3",
X"B9",
X"B3",
X"B9",
X"BB",
X"C2",
X"CE",
X"CE",
X"DA",
X"DA",
X"DA",
X"F7",
X"11",
X"1D",
X"28",
X"34",
X"3C",
X"3B",
X"40",
X"22",
X"29",
X"35",
X"33",
X"24",
X"21",
X"16",
X"06",
X"08",
X"03",
X"FA",
X"F6",
X"FA",
X"EF",
X"E8",
X"F8",
X"E4",
X"E7",
X"E8",
X"E0",
X"D7",
X"F2",
X"ED",
X"C9",
X"D2",
X"D1",
X"DE",
X"F0",
X"00",
X"F5",
X"14",
X"24",
X"1A",
X"1E",
X"17",
X"09",
X"12",
X"0E",
X"0A",
X"00",
X"F9",
X"00",
X"12",
X"1B",
X"04",
X"08",
X"F2",
X"06",
X"16",
X"09",
X"0E",
X"0C",
X"12",
X"10",
X"05",
X"00",
X"F3",
X"FE",
X"05",
X"F9",
X"00",
X"00",
X"F7",
X"EB",
X"02",
X"F0",
X"EB",
X"ED",
X"DC",
X"E3",
X"E5",
X"C8",
X"D9",
X"EA",
X"E8",
X"EE",
X"06",
X"F8",
X"FD",
X"1C",
X"22",
X"3E",
X"3C",
X"2C",
X"35",
X"18",
X"14",
X"14",
X"00",
X"00",
X"FE",
X"F8",
X"EF",
X"EF",
X"04",
X"FD",
X"EA",
X"E4",
X"E6",
X"E8",
X"EC",
X"00",
X"07",
X"12",
X"0C",
X"00",
X"35",
X"19",
X"FF",
X"00",
X"F2",
X"06",
X"E8",
X"F3",
X"CB",
X"DE",
X"FB",
X"EC",
X"05",
X"1E",
X"29",
X"31",
X"32",
X"25",
X"1D",
X"0F",
X"01",
X"FA",
X"FC",
X"01",
X"C1",
X"CA",
X"F0",
X"EB",
X"F6",
X"CF",
X"C6",
X"E9",
X"E1",
X"E2",
X"F5",
X"F7",
X"04",
X"E2",
X"F0",
X"04",
X"EC",
X"F2",
X"F2",
X"F9",
X"00",
X"13",
X"3F",
X"14",
X"34",
X"3D",
X"32",
X"30",
X"4D",
X"2F",
X"1F",
X"31",
X"11",
X"26",
X"0D",
X"07",
X"F9",
X"EF",
X"FA",
X"F3",
X"FC",
X"E4",
X"CE",
X"D3",
X"02",
X"DB",
X"AA",
X"C2",
X"BA",
X"C7",
X"BE",
X"C6",
X"C9",
X"E1",
X"E5",
X"FC",
X"08",
X"22",
X"28",
X"32",
X"48",
X"4C",
X"3E",
X"2C",
X"2D",
X"2D",
X"1F",
X"1B",
X"11",
X"FD",
X"F4",
X"EF",
X"EC",
X"FB",
X"D7",
X"F0",
X"EE",
X"FE",
X"0B",
X"0E",
X"15",
X"10",
X"11",
X"0C",
X"08",
X"04",
X"F7",
X"15",
X"0A",
X"EB",
X"00",
X"E2",
X"BB",
X"D0",
X"22",
X"E4",
X"EB",
X"03",
X"FA",
X"00",
X"F1",
X"ED",
X"DD",
X"D9",
X"D8",
X"DC",
X"CF",
X"E8",
X"E2",
X"F1",
X"10",
X"11",
X"19",
X"21",
X"33",
X"31",
X"30",
X"29",
X"3A",
X"23",
X"12",
X"13",
X"1A",
X"12",
X"07",
X"08",
X"13",
X"06",
X"12",
X"E9",
X"09",
X"0D",
X"08",
X"00",
X"F4",
X"00",
X"FB",
X"F9",
X"F7",
X"F4",
X"E9",
X"EB",
X"F5",
X"E5",
X"F1",
X"EC",
X"DA",
X"CF",
X"D6",
X"D5",
X"DF",
X"EB",
X"E1",
X"DC",
X"E2",
X"EA",
X"EB",
X"F0",
X"F3",
X"00",
X"FE",
X"07",
X"10",
X"15",
X"0B",
X"2E",
X"FF",
X"1C",
X"3C",
X"34",
X"65",
X"33",
X"38",
X"40",
X"3F",
X"35",
X"2B",
X"2F",
X"04",
X"00",
X"FD",
X"E5",
X"DC",
X"F0",
X"FB",
X"F8",
X"EC",
X"E1",
X"DA",
X"D8",
X"DC",
X"FC",
X"EF",
X"F1",
X"E1",
X"CD",
X"D3",
X"E7",
X"EC",
X"DA",
X"DD",
X"E5",
X"DE",
X"C9",
X"C4",
X"C7",
X"CA",
X"C6",
X"E7",
X"04",
X"1B",
X"30",
X"47",
X"46",
X"60",
X"5F",
X"2D",
X"4F",
X"4D",
X"2D",
X"11",
X"19",
X"0E",
X"0A",
X"1B",
X"F3",
X"06",
X"E2",
X"F7",
X"E2",
X"DB",
X"DC",
X"DE",
X"FD",
X"F9",
X"08",
X"DC",
X"11",
X"13",
X"2A",
X"12",
X"0C",
X"00",
X"FD",
X"13",
X"06",
X"F8",
X"F8",
X"FA",
X"DC",
X"DE",
X"EA",
X"D8",
X"E5",
X"E2",
X"DC",
X"D6",
X"D8",
X"B2",
X"DD",
X"EA",
X"D5",
X"12",
X"0F",
X"2C",
X"11",
X"14",
X"00",
X"05",
X"EF",
X"04",
X"0F",
X"06",
X"18",
X"1F",
X"2B",
X"33",
X"33",
X"3A",
X"4E",
X"36",
X"2B",
X"1F",
X"25",
X"16",
X"13",
X"00",
X"00",
X"EF",
X"D3",
X"DD",
X"D7",
X"DD",
X"D7",
X"D5",
X"DF",
X"DC",
X"DB",
X"D5",
X"D1",
X"EE",
X"FE",
X"E4",
X"DD",
X"02",
X"FB",
X"12",
X"F9",
X"EE",
X"13",
X"29",
X"33",
X"23",
X"29",
X"29",
X"22",
X"F7",
X"1D",
X"F5",
X"F7",
X"F2",
X"1C",
X"E5",
X"F8",
X"03",
X"DA",
X"0A",
X"F0",
X"03",
X"F3",
X"F5",
X"EE",
X"EE",
X"E8",
X"EF",
X"F0",
X"FA",
X"00",
X"09",
X"FE",
X"0B",
X"FB",
X"08",
X"12",
X"F5",
X"13",
X"20",
X"2C",
X"FE",
X"03",
X"42",
X"0E",
X"09",
X"1D",
X"01",
X"09",
X"00",
X"F8",
X"23",
X"EF",
X"FB",
X"DC",
X"BF",
X"D5",
X"EE",
X"DE",
X"E8",
X"EE",
X"E2",
X"EE",
X"F1",
X"33",
X"00",
X"15",
X"02",
X"12",
X"1D",
X"04",
X"10",
X"0C",
X"12",
X"26",
X"FD",
X"DC",
X"F0",
X"11",
X"E8",
X"E4",
X"1F",
X"F5",
X"E2",
X"09",
X"16",
X"E3",
X"F7",
X"F5",
X"F4",
X"00",
X"F7",
X"DA",
X"F5",
X"E6",
X"06",
X"E7",
X"E3",
X"05",
X"E3",
X"07",
X"00",
X"1B",
X"29",
X"22",
X"24",
X"30",
X"2B",
X"2A",
X"22",
X"21",
X"1F",
X"07",
X"1D",
X"FA",
X"E4",
X"F5",
X"FA",
X"D8",
X"D9",
X"EF",
X"E3",
X"EE",
X"ED",
X"E9",
X"04",
X"E0",
X"00",
X"FB",
X"E3",
X"00",
X"0B",
X"10",
X"F9",
X"02",
X"0B",
X"17",
X"E7",
X"00",
X"EC",
X"FB",
X"09",
X"DC",
X"FC",
X"FA",
X"04",
X"03",
X"0B",
X"05",
X"14",
X"0A",
X"EE",
X"19",
X"10",
X"FF",
X"EF",
X"DA",
X"FB",
X"F0",
X"04",
X"01",
X"16",
X"32",
X"2F",
X"36",
X"29",
X"21",
X"11",
X"00",
X"EE",
X"EB",
X"EA",
X"EA",
X"F3",
X"F2",
X"FC",
X"0E",
X"0D",
X"FF",
X"EE",
X"F4",
X"FD",
X"03",
X"DF",
X"FE",
X"F7",
X"DF",
X"F7",
X"D4",
X"C9",
X"F4",
X"E4",
X"EB",
X"FF",
X"18",
X"08",
X"F5",
X"FD",
X"F8",
X"F4",
X"FC",
X"1A",
X"0C",
X"06",
X"17",
X"0B",
X"0E",
X"24",
X"2B",
X"35",
X"30",
X"44",
X"37",
X"1F",
X"19",
X"1F",
X"24",
X"CD",
X"C7",
X"D4",
X"C6",
X"C8",
X"C3",
X"C3",
X"D6",
X"DB",
X"D7",
X"E7",
X"FB",
X"02",
X"03",
X"16",
X"2E",
X"36",
X"1A",
X"22",
X"29",
X"11",
X"0C",
X"08",
X"05",
X"E8",
X"FE",
X"01",
X"F7",
X"F3",
X"EC",
X"DC",
X"E2",
X"E0",
X"F3",
X"FA",
X"F4",
X"F9",
X"15",
X"FC",
X"F7",
X"2C",
X"2C",
X"2D",
X"3D",
X"22",
X"1C",
X"0C",
X"00",
X"F9",
X"00",
X"ED",
X"E5",
X"D7",
X"F0",
X"06",
X"BF",
X"F0",
X"E4",
X"F8",
X"F6",
X"F2",
X"F0",
X"EC",
X"E6",
X"E0",
X"D4",
X"E3",
X"EB",
X"BE",
X"ED",
X"FA",
X"06",
X"0D",
X"26",
X"1C",
X"3C",
X"45",
X"23",
X"40",
X"41",
X"4A",
X"40",
X"46",
X"31",
X"23",
X"12",
X"14",
X"F5",
X"0C",
X"13",
X"E4",
X"F7",
X"D0",
X"CD",
X"F2",
X"C6",
X"C9",
X"D2",
X"C9",
X"E2",
X"DD",
X"E6",
X"FA",
X"D0",
X"EA",
X"D0",
X"FA",
X"F7",
X"E8",
X"FA",
X"00",
X"1A",
X"0B",
X"00",
X"03",
X"F1",
X"FE",
X"15",
X"03",
X"F4",
X"0F",
X"17",
X"03",
X"15",
X"19",
X"34",
X"15",
X"21",
X"29",
X"34",
X"19",
X"01",
X"16",
X"0C",
X"0B",
X"EE",
X"E8",
X"00",
X"FF",
X"FE",
X"F9",
X"F2",
X"DD",
X"E3",
X"E7",
X"E2",
X"F0",
X"06",
X"D0",
X"13",
X"14",
X"E1",
X"00",
X"F9",
X"02",
X"15",
X"02",
X"FB",
X"00",
X"04",
X"2B",
X"F1",
X"12",
X"F7",
X"FD",
X"0C",
X"F0",
X"28",
X"0C",
X"F0",
X"FF",
X"02",
X"07",
X"E9",
X"22",
X"08",
X"CA",
X"00",
X"F2",
X"FC",
X"04",
X"FE",
X"E4",
X"F7",
X"C1",
X"00",
X"EA",
X"BB",
X"0A",
X"07",
X"0D",
X"FF",
X"16",
X"1A",
X"1D",
X"05",
X"1F",
X"F1",
X"FC",
X"11",
X"08",
X"0B",
X"05",
X"00",
X"14",
X"20",
X"14",
X"09",
X"10",
X"0C",
X"0D",
X"FA",
X"F2",
X"00",
X"03",
X"E0",
X"EA",
X"00",
X"FE",
X"FB",
X"F8",
X"FC",
X"02",
X"04",
X"07",
X"FB",
X"01",
X"FF",
X"E8",
X"EA",
X"E7",
X"E3",
X"EF",
X"FB",
X"DF",
X"F8",
X"D8",
X"05",
X"17",
X"02",
X"EC",
X"00",
X"0B",
X"EF",
X"22",
X"44",
X"FC",
X"27",
X"1C",
X"27",
X"12",
X"2B",
X"FA",
X"FD",
X"04",
X"0E",
X"F2",
X"F1",
X"09",
X"19",
X"FF",
X"FC",
X"F6",
X"ED",
X"FC",
X"EF",
X"10",
X"02",
X"F1",
X"11",
X"FC",
X"B8",
X"E1",
X"DE",
X"D3",
X"CB",
X"D7",
X"00",
X"EA",
X"EB",
X"ED",
X"E8",
X"03",
X"03",
X"12",
X"05",
X"21",
X"12",
X"1F",
X"03",
X"16",
X"17",
X"0C",
X"2A",
X"09",
X"23",
X"2E",
X"00",
X"24",
X"2D",
X"1C",
X"FA",
X"2D",
X"FC",
X"F5",
X"FA",
X"FC",
X"FC",
X"FF",
X"15",
X"FB",
X"F0",
X"EB",
X"E3",
X"E6",
X"E3",
X"F9",
X"EF",
X"B6",
X"D7",
X"F6",
X"35",
X"09",
X"E5",
X"11",
X"F0",
X"F5",
X"EB",
X"E6",
X"00",
X"E8",
X"00",
X"24",
X"E6",
X"DF",
X"02",
X"F5",
X"FF",
X"0F",
X"1C",
X"FB",
X"00",
X"02",
X"20",
X"00",
X"F5",
X"0A",
X"F7",
X"13",
X"FB",
X"F4",
X"0C",
X"08",
X"20",
X"F6",
X"E2",
X"14",
X"FE",
X"00",
X"17",
X"2E",
X"11",
X"0B",
X"14",
X"FA",
X"04",
X"03",
X"F1",
X"01",
X"F0",
X"EF",
X"F5",
X"F5",
X"FB",
X"00",
X"0B",
X"0A",
X"12",
X"17",
X"15",
X"1F",
X"1F",
X"04",
X"0B",
X"05",
X"06",
X"F9",
X"F4",
X"F0",
X"E3",
X"E6",
X"B3",
X"D1",
X"E8",
X"E8",
X"F2",
X"FC",
X"F1",
X"E2",
X"E2",
X"DB",
X"D4",
X"D9",
X"DE",
X"DF",
X"04",
X"36",
X"2A",
X"1F",
X"24",
X"19",
X"2B",
X"42",
X"3C",
X"4C",
X"46",
X"25",
X"17",
X"24",
X"44",
X"E4",
X"C6",
X"EA",
X"E0",
X"B8",
X"CF",
X"CD",
X"E0",
X"E6",
X"EC",
X"ED",
X"00",
X"00",
X"0E",
X"2A",
X"1C",
X"13",
X"32",
X"29",
X"16",
X"0F",
X"00",
X"CE",
X"F8",
X"D1",
X"EB",
X"E6",
X"C0",
X"EB",
X"E5",
X"FB",
X"F7",
X"00",
X"03",
X"FB",
X"FF",
X"03",
X"05",
X"00",
X"01",
X"0C",
X"13",
X"13",
X"44",
X"03",
X"F5",
X"20",
X"0F",
X"38",
X"02",
X"19",
X"FE",
X"02",
X"FB",
X"F8",
X"0B",
X"F1",
X"EC",
X"C2",
X"A4",
X"CB",
X"F3",
X"E7",
X"E4",
X"04",
X"01",
X"14",
X"15",
X"06",
X"E0",
X"E9",
X"FB",
X"FD",
X"05",
X"0F",
X"0E",
X"24",
X"15",
X"06",
X"25",
X"20",
X"EE",
X"0F",
X"16",
X"0A",
X"15",
X"22",
X"3D",
X"20",
X"16",
X"EC",
X"0E",
X"32",
X"FC",
X"12",
X"F7",
X"12",
X"FB",
X"F4",
X"BF",
X"C1",
X"CE",
X"BB",
X"B1",
X"D0",
X"D4",
X"D7",
X"D6",
X"E2",
X"E7",
X"12",
X"25",
X"F4",
X"03",
X"F5",
X"07",
X"1E",
X"32",
X"62",
X"2B",
X"1E",
X"27",
X"28",
X"18",
X"17",
X"05",
X"EF",
X"0B",
X"05",
X"D6",
X"BD",
X"F5",
X"F5",
X"28",
X"EC",
X"FB",
X"F7",
X"F7",
X"F5",
X"DD",
X"E8",
X"F3",
X"F2",
X"C4",
X"E1",
X"FA",
X"F7",
X"F5",
X"03",
X"33",
X"0D",
X"01",
X"43",
X"44",
X"FF",
X"22",
X"15",
X"0A",
X"1E",
X"38",
X"EE",
X"F3",
X"0D",
X"CC",
X"21",
X"08",
X"11",
X"F8",
X"D1",
X"00",
X"F1",
X"03",
X"15",
X"15",
X"DB",
X"CC",
X"F3",
X"C4",
X"C2",
X"1C",
X"EC",
X"CA",
X"F6",
X"00",
X"EE",
X"EE",
X"F9",
X"F9",
X"B5",
X"FD",
X"EE",
X"F6",
X"0E",
X"22",
X"35",
X"22",
X"23",
X"21",
X"22",
X"1B",
X"20",
X"1B",
X"24",
X"19",
X"1C",
X"18",
X"3D",
X"14",
X"0C",
X"00",
X"0C",
X"04",
X"E5",
X"FF",
X"E3",
X"08",
X"08",
X"1C",
X"02",
X"DF",
X"DE",
X"C4",
X"B3",
X"B6",
X"BA",
X"C0",
X"CC",
X"ED",
X"E7",
X"00",
X"0D",
X"11",
X"2A",
X"1A",
X"10",
X"18",
X"0F",
X"1D",
X"15",
X"0C",
X"FA",
X"FB",
X"F3",
X"CC",
X"FB",
X"D7",
X"F9",
X"E2",
X"EE",
X"F1",
X"09",
X"0C",
X"FF",
X"23",
X"25",
X"04",
X"31",
X"1E",
X"2F",
X"28",
X"4A",
X"30",
X"43",
X"48",
X"00",
X"1E",
X"0D",
X"28",
X"FE",
X"DF",
X"0B",
X"D9",
X"FF",
X"E8",
X"CB",
X"E9",
X"9B",
X"B5",
X"AB",
X"C6",
X"BF",
X"C8",
X"C5",
X"FD",
X"FF",
X"E9",
X"00",
X"0C",
X"F5",
X"ED",
X"06",
X"00",
X"33",
X"13",
X"0F",
X"2E",
X"28",
X"1D",
X"07",
X"13",
X"52",
X"3A",
X"03",
X"19",
X"EF",
X"00",
X"27",
X"1A",
X"ED",
X"30",
X"12",
X"FB",
X"DF",
X"F4",
X"F3",
X"C8",
X"D8",
X"DC",
X"FE",
X"FC",
X"D1",
X"02",
X"04",
X"D4",
X"02",
X"04",
X"1A",
X"0A",
X"EF",
X"11",
X"F5",
X"F3",
X"2D",
X"E8",
X"C5",
X"D4",
X"FA",
X"03",
X"08",
X"01",
X"36",
X"06",
X"18",
X"26",
X"EF",
X"00",
X"26",
X"D6",
X"25",
X"F6",
X"08",
X"00",
X"16",
X"02",
X"30",
X"05",
X"E6",
X"2B",
X"36",
X"D9",
X"F2",
X"EE",
X"F7",
X"EC",
X"E8",
X"00",
X"CA",
X"FB",
X"F8",
X"C0",
X"B7",
X"C8",
X"E7",
X"E3",
X"E7",
X"1A",
X"FA",
X"16",
X"15",
X"22",
X"13",
X"23",
X"0B",
X"0B",
X"12",
X"05",
X"FF",
X"FA",
X"0D",
X"18",
X"F6",
X"20",
X"14",
X"16",
X"0D",
X"20",
X"F5",
X"0C",
X"0F",
X"0E",
X"00",
X"FC",
X"F3",
X"1A",
X"D6",
X"00",
X"FF",
X"33",
X"00",
X"FB",
X"0E",
X"0C",
X"D3",
X"0F",
X"DA",
X"DE",
X"E0",
X"CA",
X"DE",
X"DD",
X"11",
X"F4",
X"D4",
X"BA",
X"02",
X"FE",
X"14",
X"FE",
X"21",
X"0C",
X"13",
X"20",
X"0F",
X"24",
X"3A",
X"F6",
X"2A",
X"F1",
X"3B",
X"0B",
X"EE",
X"07",
X"04",
X"16",
X"F6",
X"FA",
X"04",
X"15",
X"DF",
X"F0",
X"FD",
X"DE",
X"D3",
X"D1",
X"E3",
X"C1",
X"BA",
X"EA",
X"F7",
X"12",
X"28",
X"0B",
X"E7",
X"FC",
X"00",
X"EB",
X"E7",
X"10",
X"F6",
X"DC",
X"21",
X"34",
X"EB",
X"1F",
X"36",
X"5C",
X"06",
X"00",
X"36",
X"1D",
X"2C",
X"0B",
X"22",
X"19",
X"14",
X"0D",
X"FD",
X"04",
X"F8",
X"EC",
X"CC",
X"FE",
X"DB",
X"E7",
X"FB",
X"FE",
X"03",
X"0B",
X"09",
X"DF",
X"DB",
X"F0",
X"FC",
X"45",
X"15",
X"D2",
X"09",
X"09",
X"07",
X"D2",
X"F0",
X"E8",
X"C3",
X"E2",
X"D1",
X"C3",
X"DE",
X"E3",
X"D6",
X"DB",
X"FE",
X"F0",
X"30",
X"22",
X"0B",
X"16",
X"4F",
X"3A",
X"FD",
X"34",
X"4C",
X"4E",
X"02",
X"FC",
X"FC",
X"D4",
X"23",
X"D9",
X"F2",
X"00",
X"F9",
X"00",
X"EA",
X"EB",
X"09",
X"D3",
X"D0",
X"1D",
X"0B",
X"C2",
X"F0",
X"16",
X"34",
X"1B",
X"11",
X"20",
X"31",
X"20",
X"10",
X"00",
X"F6",
X"D4",
X"C8",
X"E5",
X"DC",
X"F9",
X"F0",
X"15",
X"FB",
X"F7",
X"E8",
X"12",
X"DA",
X"E4",
X"04",
X"1A",
X"37",
X"12",
X"34",
X"29",
X"1E",
X"1E",
X"25",
X"19",
X"1C",
X"13",
X"06",
X"FE",
X"F1",
X"FC",
X"F5",
X"D0",
X"C8",
X"E7",
X"0B",
X"D4",
X"BE",
X"EA",
X"E0",
X"E2",
X"DD",
X"E7",
X"D1",
X"ED",
X"F3",
X"A4",
X"E8",
X"C8",
X"D8",
X"16",
X"40",
X"2A",
X"F9",
X"3C",
X"13",
X"2B",
X"21",
X"41",
X"55",
X"35",
X"52",
X"3F",
X"FF",
X"2E",
X"F7",
X"0C",
X"2E",
X"FE",
X"0F",
X"E6",
X"F7",
X"C2",
X"B0",
X"C5",
X"D8",
X"E5",
X"EF",
X"FB",
X"EE",
X"FB",
X"E6",
X"E2",
X"E1",
X"F6",
X"F5",
X"0D",
X"1E",
X"26",
X"19",
X"49",
X"10",
X"2F",
X"34",
X"46",
X"0E",
X"F2",
X"1A",
X"DE",
X"FD",
X"ED",
X"0D",
X"D5",
X"DD",
X"E0",
X"BD",
X"C6",
X"C2",
X"BA",
X"D2",
X"F6",
X"BF",
X"C3",
X"F5",
X"02",
X"0C",
X"41",
X"05",
X"1F",
X"26",
X"24",
X"2F",
X"19",
X"FF",
X"27",
X"FE",
X"F0",
X"44",
X"38",
X"30",
X"E8",
X"35",
X"15",
X"F5",
X"09",
X"FC",
X"01",
X"E2",
X"0A",
X"FA",
X"04",
X"F9",
X"B8",
X"F3",
X"CC",
X"F3",
X"0B",
X"07",
X"24",
X"15",
X"20",
X"00",
X"2F",
X"F9",
X"D6",
X"DE",
X"A2",
X"CD",
X"CB",
X"D9",
X"06",
X"FF",
X"03",
X"DC",
X"E5",
X"2D",
X"E1",
X"20",
X"1F",
X"4E",
X"EE",
X"F8",
X"35",
X"37",
X"1E",
X"F0",
X"F9",
X"32",
X"50",
X"00",
X"FD",
X"20",
X"08",
X"C9",
X"43",
X"EE",
X"19",
X"F2",
X"E4",
X"F3",
X"0D",
X"07",
X"C5",
X"13",
X"C1",
X"C1",
X"F9",
X"D0",
X"AA",
X"F7",
X"11",
X"08",
X"F2",
X"BF",
X"DC",
X"1C",
X"DD",
X"F2",
X"26",
X"0C",
X"DC",
X"F9",
X"EF",
X"08",
X"0F",
X"E4",
X"3E",
X"21",
X"53",
X"34",
X"2A",
X"28",
X"2B",
X"1D",
X"37",
X"25",
X"19",
X"E3",
X"DD",
X"FB",
X"EE",
X"12",
X"B5",
X"E0",
X"C4",
X"FB",
X"3C",
X"E8",
X"E8",
X"3A",
X"EE",
X"0F",
X"15",
X"05",
X"ED",
X"15",
X"06",
X"C3",
X"E3",
X"D8",
X"E0",
X"D9",
X"F5",
X"D5",
X"20",
X"FC",
X"DF",
X"3E",
X"DB",
X"CF",
X"17",
X"19",
X"FF",
X"DD",
X"0E",
X"14",
X"20",
X"E7",
X"05",
X"20",
X"C4",
X"CB",
X"0C",
X"23",
X"1A",
X"25",
X"56",
X"1A",
X"29",
X"04",
X"00",
X"06",
X"E9",
X"E2",
X"EA",
X"0C",
X"16",
X"2A",
X"15",
X"F3",
X"15",
X"0C",
X"DB",
X"D4",
X"12",
X"35",
X"D4",
X"AD",
X"C7",
X"25",
X"E6",
X"E1",
X"0C",
X"0A",
X"0F",
X"E1",
X"C8",
X"F3",
X"FA",
X"E3",
X"E5",
X"05",
X"0D",
X"23",
X"20",
X"1B",
X"2F",
X"2B",
X"EA",
X"D1",
X"09",
X"0C",
X"F8",
X"03",
X"17",
X"14",
X"0A",
X"1C",
X"2B",
X"DD",
X"BB",
X"E3",
X"E1",
X"DA",
X"10",
X"FF",
X"E6",
X"EC",
X"04",
X"15",
X"44",
X"49",
X"41",
X"37",
X"2C",
X"0C",
X"01",
X"E8",
X"E8",
X"D7",
X"E7",
X"F0",
X"EA",
X"EC",
X"BD",
X"D6",
X"F1",
X"F2",
X"2A",
X"39",
X"14",
X"13",
X"D3",
X"F2",
X"00",
X"21",
X"13",
X"F0",
X"F4",
X"E2",
X"D4",
X"DF",
X"DE",
X"FB",
X"D2",
X"F9",
X"0F",
X"C8",
X"E2",
X"F8",
X"F7",
X"03",
X"05",
X"10",
X"0B",
X"07",
X"0D",
X"1A",
X"2B",
X"14",
X"1C",
X"1E",
X"01",
X"06",
X"0F",
X"14",
X"1F",
X"54",
X"2E",
X"39",
X"46",
X"06",
X"E6",
X"E4",
X"29",
X"27",
X"F1",
X"11",
X"24",
X"E6",
X"FC",
X"DA",
X"FC",
X"BC",
X"C5",
X"05",
X"AB",
X"8B",
X"94",
X"E4",
X"DF",
X"C3",
X"F7",
X"EE",
X"15",
X"10",
X"0B",
X"12",
X"0C",
X"E5",
X"EF",
X"E7",
X"04",
X"EA",
X"D4",
X"34",
X"F2",
X"19",
X"00",
X"26",
X"19",
X"12",
X"39",
X"41",
X"09",
X"F5",
X"26",
X"52",
X"30",
X"22",
X"24",
X"E0",
X"04",
X"25",
X"33",
X"1A",
X"D5",
X"EA",
X"18",
X"00",
X"16",
X"F9",
X"FF",
X"CC",
X"C8",
X"BC",
X"CF",
X"E3",
X"DC",
X"E0",
X"B7",
X"E3",
X"11",
X"0A",
X"1F",
X"EA",
X"F5",
X"20",
X"0D",
X"BF",
X"F5",
X"F6",
X"ED",
X"17",
X"0B",
X"00",
X"18",
X"42",
X"FA",
X"D7",
X"EA",
X"DB",
X"00",
X"07",
X"11",
X"1D",
X"13",
X"4A",
X"2B",
X"02",
X"27",
X"32",
X"FD",
X"03",
X"06",
X"3F",
X"D5",
X"13",
X"0A",
X"A1",
X"04",
X"D6",
X"05",
X"19",
X"25",
X"00",
X"CD",
X"EE",
X"E3",
X"DF",
X"FC",
X"E1",
X"FC",
X"CC",
X"C2",
X"38",
X"E2",
X"BE",
X"34",
X"1C",
X"C8",
X"1B",
X"00",
X"FA",
X"F6",
X"33",
X"CA",
X"03",
X"12",
X"DF",
X"31",
X"1A",
X"03",
X"20",
X"1B",
X"1A",
X"F7",
X"EB",
X"10",
X"21",
X"23",
X"26",
X"19",
X"0E",
X"23",
X"DF",
X"EB",
X"D6",
X"FE",
X"F5",
X"D6",
X"EF",
X"FD",
X"EF",
X"FB",
X"09",
X"04",
X"00",
X"25",
X"16",
X"FA",
X"EB",
X"DF",
X"FB",
X"0D",
X"18",
X"54",
X"3A",
X"E7",
X"14",
X"0F",
X"F9",
X"D0",
X"B5",
X"EC",
X"DB",
X"30",
X"05",
X"A4",
X"1B",
X"08",
X"CF",
X"E5",
X"F4",
X"BB",
X"D5",
X"EC",
X"00",
X"2D",
X"4F",
X"F5",
X"D6",
X"F8",
X"FE",
X"00",
X"E4",
X"09",
X"F3",
X"13",
X"05",
X"31",
X"00",
X"31",
X"38",
X"13",
X"4E",
X"12",
X"D1",
X"08",
X"07",
X"EA",
X"1B",
X"FF",
X"FE",
X"11",
X"1F",
X"2B",
X"27",
X"09",
X"0F",
X"09",
X"31",
X"1B",
X"D3",
X"F3",
X"04",
X"F4",
X"D9",
X"BF",
X"BB",
X"C6",
X"CE",
X"AD",
X"A3",
X"CB",
X"D7",
X"E3",
X"00",
X"24",
X"29",
X"EA",
X"FC",
X"0C",
X"1C",
X"24",
X"FC",
X"05",
X"0A",
X"25",
X"FD",
X"12",
X"3D",
X"3F",
X"01",
X"00",
X"15",
X"47",
X"30",
X"1B",
X"0E",
X"EF",
X"06",
X"E7",
X"F0",
X"0F",
X"EC",
X"CF",
X"CC",
X"F0",
X"F3",
X"E2",
X"DF",
X"DA",
X"FE",
X"05",
X"0C",
X"FA",
X"14",
X"10",
X"FA",
X"EC",
X"FD",
X"00",
X"03",
X"04",
X"00",
X"2A",
X"14",
X"DF",
X"20",
X"08",
X"FF",
X"20",
X"34",
X"0B",
X"FD",
X"17",
X"0B",
X"13",
X"18",
X"1C",
X"F1",
X"0B",
X"C1",
X"A8",
X"E0",
X"D2",
X"F1",
X"D4",
X"DC",
X"CD",
X"D9",
X"DF",
X"09",
X"11",
X"E7",
X"F9",
X"ED",
X"08",
X"E4",
X"22",
X"40",
X"52",
X"0A",
X"00",
X"27",
X"40",
X"56",
X"41",
X"24",
X"FC",
X"18",
X"E9",
X"E2",
X"28",
X"03",
X"CB",
X"07",
X"F4",
X"02",
X"EF",
X"FC",
X"07",
X"F2",
X"B9",
X"DE",
X"C1",
X"F9",
X"03",
X"08",
X"F7",
X"E9",
X"BF",
X"DF",
X"F9",
X"B8",
X"06",
X"04",
X"F3",
X"13",
X"2C",
X"1E",
X"17",
X"1A",
X"FB",
X"D3",
X"F0",
X"D7",
X"00",
X"12",
X"43",
X"32",
X"FC",
X"19",
X"31",
X"05",
X"16",
X"08",
X"20",
X"F6",
X"8E",
X"CF",
X"F2",
X"00",
X"28",
X"16",
X"F9",
X"0C",
X"0B",
X"14",
X"01",
X"ED",
X"09",
X"17",
X"EE",
X"1C",
X"53",
X"09",
X"0D",
X"1B",
X"08",
X"15",
X"0A",
X"FA",
X"F1",
X"DE",
X"EB",
X"11",
X"01",
X"97",
X"A3",
X"DF",
X"ED",
X"04",
X"0E",
X"19",
X"14",
X"08",
X"FD",
X"0B",
X"00",
X"CC",
X"E3",
X"C5",
X"CB",
X"02",
X"E4",
X"E4",
X"11",
X"09",
X"FC",
X"1E",
X"0F",
X"1F",
X"1B",
X"25",
X"16",
X"30",
X"20",
X"FD",
X"1E",
X"11",
X"E5",
X"12",
X"40",
X"EC",
X"09",
X"2F",
X"F3",
X"36",
X"3A",
X"E1",
X"04",
X"F8",
X"DF",
X"C3",
X"05",
X"DA",
X"D7",
X"00",
X"D6",
X"F8",
X"F8",
X"E4",
X"EA",
X"B1",
X"DB",
X"CD",
X"DB",
X"F2",
X"18",
X"E2",
X"F7",
X"0C",
X"11",
X"10",
X"31",
X"2E",
X"00",
X"16",
X"35",
X"4A",
X"29",
X"E4",
X"11",
X"62",
X"F9",
X"FE",
X"03",
X"19",
X"19",
X"44",
X"15",
X"FC",
X"FF",
X"02",
X"EE",
X"D8",
X"D5",
X"96",
X"BB",
X"0C",
X"F9",
X"E8",
X"B8",
X"DD",
X"EF",
X"18",
X"03",
X"2A",
X"22",
X"D1",
X"06",
X"F2",
X"F6",
X"FC",
X"F9",
X"E9",
X"AC",
X"EA",
X"0E",
X"E4",
X"ED",
X"4A",
X"3F",
X"18",
X"FB",
X"F6",
X"64",
X"14",
X"F9",
X"33",
X"E9",
X"0E",
X"2C",
X"00",
X"F8",
X"D9",
X"F0",
X"ED",
X"13",
X"13",
X"00",
X"3D",
X"1D",
X"FD",
X"0B",
X"FD",
X"00",
X"00",
X"03",
X"0D",
X"04",
X"00",
X"FB",
X"12",
X"D8",
X"E1",
X"DB",
X"D4",	
X"D4" );
--//--------------------------------------
  begin

    if (RESET_N='0') then
      Q <= sqr_table(0);
    elsif(rising_edge(CLK)) then
      if (ENA='1') then
          Q <= sqr_table(to_integer(unsigned(ADDR)));
      end if;
    end if;
  end process;
end arch;