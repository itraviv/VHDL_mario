--------------------------------------
-- SinTable.vhd
-- Written by Saar Eliad and Itamar Raviv.
-- All rights reserved, Copyright 2017
--------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity goldSoundTable is
port(
  CLK     : in std_logic;
  RESET_N : in std_logic;
  ENA     : in std_logic;
  ADDR    : in std_logic_vector(11 downto 0);
  Q       : out std_logic_vector(7 downto 0)
);
end goldSoundTable;

architecture arch of goldSoundTable is

type table_type is array(0 to 4095) of std_logic_vector(7 downto 0);
signal sqr_table : table_type;

begin

  goldSoundTable_proc: process(RESET_N, CLK)
    constant sqr_table : table_type := (
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"02",
X"FE",
X"03",
X"DF",
X"81",
X"93",
X"88",
X"D3",
X"21",
X"10",
X"20",
X"EB",
X"93",
X"A8",
X"9E",
X"D3",
X"31",
X"25",
X"2F",
X"09",
X"AC",
X"AD",
X"A7",
X"CC",
X"31",
X"37",
X"3B",
X"25",
X"BF",
X"B4",
X"B8",
X"CB",
X"33",
X"48",
X"44",
X"3B",
X"D8",
X"B7",
X"C2",
X"C7",
X"2C",
X"55",
X"48",
X"4D",
X"F0",
X"BC",
X"CA",
X"C5",
X"21",
X"5D",
X"50",
X"59",
X"05",
X"C0",
X"D3",
X"C9",
X"17",
X"62",
X"52",
X"5D",
X"1B",
X"C6",
X"D4",
X"C9",
X"01",
X"5D",
X"54",
X"5E",
X"30",
X"CE",
X"D4",
X"CD",
X"F7",
X"58",
X"56",
X"5C",
X"40",
X"D9",
X"D3",
X"CF",
X"E6",
X"4C",
X"56",
X"56",
X"4C",
X"E7",
X"D1",
X"D3",
X"D9",
X"3C",
X"57",
X"4E",
X"51",
X"F0",
X"CA",
X"D3",
X"CF",
X"2A",
X"56",
X"49",
X"54",
X"00",
X"C6",
X"D2",
X"C5",
X"16",
X"54",
X"46",
X"53",
X"0D",
X"C3",
X"D1",
X"C1",
X"01",
X"50",
X"44",
X"53",
X"1B",
X"C3",
X"CE",
X"BE",
X"F1",
X"4A",
X"44",
X"51",
X"2B",
X"CA",
X"CC",
X"C0",
X"E0",
X"41",
X"45",
X"4C",
X"37",
X"D1",
X"C7",
X"C3",
X"D1",
X"34",
X"42",
X"40",
X"3C",
X"DB",
X"C2",
X"C6",
X"C5",
X"24",
X"42",
X"3C",
X"42",
X"E9",
X"BF",
X"C8",
X"BE",
X"15",
X"43",
X"39",
X"45",
X"F9",
X"BC",
X"C9",
X"BB",
X"04",
X"44",
X"37",
X"44",
X"04",
X"BA",
X"C7",
X"B8",
X"F4",
X"3F",
X"34",
X"41",
X"12",
X"BE",
X"C6",
X"B9",
X"E3",
X"38",
X"32",
X"3B",
X"1C",
X"C0",
X"BF",
X"B8",
X"D2",
X"2F",
X"35",
X"38",
X"28",
X"CA",
X"BB",
X"BB",
X"C5",
X"22",
X"36",
X"31",
X"2F",
X"D5",
X"B6",
X"BE",
X"BB",
X"14",
X"38",
X"2D",
X"36",
X"E3",
X"B4",
X"B8",
X"AA",
X"FE",
X"30",
X"2E",
X"39",
X"F3",
X"B4",
X"B9",
X"AC",
X"F2",
X"32",
X"30",
X"3D",
X"08",
X"B7",
X"B5",
X"A7",
X"DB",
X"2E",
X"33",
X"3E",
X"19",
X"C0",
X"B8",
X"AE",
X"CF",
X"2A",
X"35",
X"3D",
X"28",
X"CA",
X"B9",
X"B5",
X"C5",
X"23",
X"37",
X"39",
X"32",
X"D7",
X"B8",
X"B8",
X"BA",
X"15",
X"3A",
X"36",
X"3A",
X"E7",
X"B9",
X"BE",
X"B6",
X"04",
X"38",
X"31",
X"3C",
X"F6",
X"B5",
X"BB",
X"B1",
X"F6",
X"38",
X"32",
X"40",
X"09",
X"BD",
X"C1",
X"B1",
X"E4",
X"33",
X"31",
X"3F",
X"17",
X"C2",
X"BF",
X"B1",
X"D3",
X"29",
X"2C",
X"36",
X"20",
X"C7",
X"BA",
X"B0",
X"C3",
X"1D",
X"2F",
X"34",
X"2C",
X"D3",
X"BB",
X"B6",
X"BD",
X"13",
X"31",
X"31",
X"33",
X"E0",
X"BA",
X"BC",
X"B8",
X"0A",
X"37",
X"31",
X"3A",
X"EE",
X"B8",
X"BD",
X"B3",
X"FD",
X"37",
X"30",
X"3D",
X"FE",
X"BB",
X"C1",
X"B2",
X"EE",
X"34",
X"2E",
X"3C",
X"0D",
X"BE",
X"C1",
X"B2",
X"DE",
X"2F",
X"2F",
X"3B",
X"1C",
X"C6",
X"C0",
X"B4",
X"D0",
X"28",
X"32",
X"38",
X"27",
X"CE",
X"BD",
X"B7",
X"C2",
X"1B",
X"32",
X"34",
X"34",
X"DB",
X"BC",
X"BC",
X"BB",
X"11",
X"35",
X"32",
X"3A",
X"EA",
X"BE",
X"C4",
X"B9",
X"07",
X"39",
X"30",
X"3F",
X"F9",
X"C0",
X"C7",
X"B8",
X"FB",
X"38",
X"2D",
X"3F",
X"06",
X"C1",
X"C8",
X"B7",
X"EB",
X"36",
X"2E",
X"3F",
X"17",
X"C8",
X"CB",
X"BB",
X"DD",
X"2E",
X"2D",
X"3A",
X"24",
X"CF",
X"CA",
X"BF",
X"D0",
X"27",
X"2E",
X"36",
X"2F",
X"D9",
X"C9",
X"C2",
X"C5",
X"1C",
X"32",
X"33",
X"3A",
X"E7",
X"C9",
X"CA",
X"BE",
X"10",
X"34",
X"2E",
X"41",
X"F6",
X"C9",
X"D0",
X"BD",
X"05",
X"39",
X"2D",
X"42",
X"00",
X"C6",
X"D3",
X"BE",
X"FB",
X"3A",
X"2E",
X"45",
X"13",
X"CC",
X"D6",
X"C1",
X"ED",
X"3A",
X"30",
X"45",
X"23",
X"CE",
X"D4",
X"C2",
X"DF",
X"38",
X"34",
X"44",
X"32",
X"D6",
X"D1",
X"C5",
X"D1",
X"30",
X"38",
X"40",
X"3E",
X"E1",
X"CE",
X"CB",
X"C9",
X"28",
X"3D",
X"3C",
X"44",
X"EE",
X"D0",
X"D5",
X"C6",
X"19",
X"3C",
X"37",
X"49",
X"FF",
X"CE",
X"D7",
X"BF",
X"09",
X"3C",
X"31",
X"49",
X"0A",
X"CA",
X"D8",
X"BD",
X"FC",
X"3B",
X"2E",
X"46",
X"17",
X"CB",
X"DB",
X"BE",
X"EC",
X"38",
X"2E",
X"43",
X"26",
X"CF",
X"D7",
X"C1",
X"DB",
X"34",
X"2F",
X"40",
X"35",
X"D5",
X"D4",
X"C7",
X"D0",
X"2E",
X"33",
X"39",
X"3A",
X"DF",
X"D1",
X"CD",
X"C7",
X"21",
X"36",
X"33",
X"42",
X"EC",
X"CD",
X"D3",
X"BF",
X"14",
X"37",
X"2E",
X"44",
X"FA",
X"C9",
X"D7",
X"BB",
X"04",
X"39",
X"2A",
X"44",
X"07",
X"C7",
X"D9",
X"BA",
X"F7",
X"37",
X"28",
X"42",
X"17",
X"C7",
X"D9",
X"BB",
X"E6",
X"35",
X"29",
X"3E",
X"24",
X"CD",
X"D7",
X"C1",
X"D9",
X"2F",
X"2C",
X"38",
X"31",
X"D5",
X"D5",
X"C7",
X"CE",
X"27",
X"31",
X"33",
X"3C",
X"E0",
X"D2",
X"CF",
X"C5",
X"1B",
X"36",
X"2B",
X"43",
X"EB",
X"CD",
X"D3",
X"C2",
X"0F",
X"3A",
X"28",
X"47",
X"FC",
X"CC",
X"D6",
X"BE",
X"FD",
X"3C",
X"26",
X"48",
X"08",
X"C9",
X"D5",
X"BF",
X"EE",
X"3E",
X"25",
X"45",
X"16",
X"CD",
X"D4",
X"C4",
X"E0",
X"39",
X"26",
X"40",
X"23",
X"D2",
X"D0",
X"C9",
X"D2",
X"34",
X"2A",
X"39",
X"2F",
X"DA",
X"CB",
X"D1",
X"C6",
X"2B",
X"30",
X"37",
X"36",
X"EB",
X"C7",
X"D7",
X"BD",
X"23",
X"2F",
X"3C",
X"13",
X"C6",
X"CC",
X"F9",
X"30",
X"40",
X"13",
X"C7",
X"D4",
X"E3",
X"3D",
X"3D",
X"19",
X"D3",
X"CB",
X"DA",
X"3D",
X"31",
X"22",
X"D9",
X"C8",
X"E5",
X"3B",
X"2B",
X"2E",
X"CA",
X"C7",
X"E4",
X"31",
X"3A",
X"35",
X"C8",
X"CC",
X"D0",
X"26",
X"42",
X"35",
X"E0",
X"D6",
X"C2",
X"21",
X"32",
X"2D",
X"ED",
X"D3",
X"CF",
X"28",
X"2A",
X"30",
X"E7",
X"C3",
X"D4",
X"21",
X"36",
X"3F",
X"EB",
X"C0",
X"CC",
X"08",
X"3B",
X"40",
X"F8",
X"D3",
X"C9",
X"00",
X"38",
X"2E",
X"00",
X"D3",
X"CC",
X"08",
X"3C",
X"2C",
X"08",
X"BD",
X"CA",
X"00",
X"3D",
X"3C",
X"16",
X"C0",
X"CD",
X"E9",
X"33",
X"38",
X"1B",
X"CD",
X"D8",
X"E3",
X"39",
X"2C",
X"16",
X"CB",
X"D4",
X"E5",
X"42",
X"2D",
X"23",
X"C8",
X"C6",
X"D7",
X"39",
X"34",
X"37",
X"CF",
X"C9",
X"CC",
X"24",
X"2D",
X"37",
X"DA",
X"DA",
X"D0",
X"23",
X"29",
X"2C",
X"D7",
X"D7",
X"D3",
X"2C",
X"33",
X"2E",
X"DA",
X"C7",
X"C6",
X"23",
X"39",
X"3D",
X"EE",
X"C8",
X"C2",
X"0F",
X"2E",
X"3A",
X"FA",
X"D1",
X"CE",
X"09",
X"2C",
X"32",
X"F6",
X"CA",
X"D0",
X"06",
X"3B",
X"36",
X"FD",
X"C3",
X"C3",
X"F7",
X"3E",
X"39",
X"12",
X"CB",
X"C4",
X"EB",
X"32",
X"2E",
X"1D",
X"CF",
X"D1",
X"EB",
X"2F",
X"29",
X"1B",
X"C5",
X"D5",
X"E5",
X"37",
X"32",
X"1E",
X"C3",
X"CF",
X"D3",
X"39",
X"32",
X"2C",
X"D2",
X"CE",
X"CB",
X"31",
X"25",
X"32",
X"D9",
X"D3",
X"D3",
X"2A",
X"20",
X"30",
X"D2",
X"D3",
X"D5",
X"27",
X"2D",
X"32",
X"D1",
X"D0",
X"C8",
X"1F",
X"35",
X"34",
X"E6",
X"CB",
X"BE",
X"15",
X"2F",
X"39",
X"F5",
X"CB",
X"C4",
X"09",
X"27",
X"36",
X"FA",
X"CC",
X"CF",
X"02",
X"2F",
X"2F",
X"F8",
X"CB",
X"CE",
X"00",
X"39",
X"27",
X"00",
X"C6",
X"CE",
X"FF",
X"3A",
X"29",
X"07",
X"BC",
X"CE",
X"F7",
X"3A",
X"31",
X"10",
X"BC",
X"CF",
X"E5",
X"38",
X"2F",
X"17",
X"C8",
X"D3",
X"DE",
X"35",
X"24",
X"18",
X"CE",
X"D1",
X"E1",
X"35",
X"20",
X"1D",
X"C8",
X"CE",
X"E1",
X"30",
X"28",
X"24",
X"C7",
X"D0",
X"D9",
X"29",
X"2D",
X"25",
X"D2",
X"D3",
X"D0",
X"24",
X"28",
X"24",
X"DD",
X"D4",
X"D3",
X"25",
X"26",
X"23",
X"DE",
X"CC",
X"D5",
X"20",
X"2C",
X"2D",
X"E5",
X"C7",
X"CF",
X"0E",
X"2F",
X"31",
X"F1",
X"CF",
X"CF",
X"02",
X"2C",
X"27",
X"FA",
X"D7",
X"DA",
X"07",
X"32",
X"21",
X"FD",
X"CB",
X"D5",
X"03",
X"36",
X"27",
X"07",
X"C5",
X"D3",
X"F6",
X"31",
X"28",
X"0F",
X"CB",
X"DB",
X"EB",
X"2E",
X"21",
X"0D",
X"CB",
X"DD",
X"EA",
X"35",
X"1E",
X"10",
X"C5",
X"D4",
X"E3",
X"38",
X"23",
X"1F",
X"C8",
X"D0",
X"D8",
X"2D",
X"22",
X"26",
X"CE",
X"D8",
X"D6",
X"27",
X"1E",
X"21",
X"D1",
X"DA",
X"D7",
X"2B",
X"22",
X"20",
X"CF",
X"D1",
X"D1",
X"28",
X"28",
X"2A",
X"DA",
X"CD",
X"CC",
X"19",
X"25",
X"2B",
X"E6",
X"D1",
X"D4",
X"12",
X"25",
X"23",
X"E6",
X"CD",
X"D7",
X"11",
X"31",
X"24",
X"EC",
X"C4",
X"CF",
X"05",
X"37",
X"28",
X"FE",
X"C6",
X"CE",
X"F9",
X"2E",
X"22",
X"07",
X"CB",
X"DD",
X"F6",
X"2E",
X"18",
X"04",
X"C1",
X"E0",
X"F6",
X"3D",
X"20",
X"09",
X"B9",
X"D4",
X"E6",
X"40",
X"26",
X"1D",
X"C3",
X"D2",
X"D8",
X"32",
X"1C",
X"25",
X"CC",
X"E0",
X"DC",
X"30",
X"17",
X"1C",
X"C4",
X"DE",
X"DE",
X"36",
X"23",
X"23",
X"C6",
X"D3",
X"CF",
X"2E",
X"28",
X"2D",
X"D9",
X"D5",
X"CB",
X"1F",
X"1D",
X"29",
X"E3",
X"DB",
X"D8",
X"1B",
X"1F",
X"21",
X"E1",
X"D5",
X"DA",
X"19",
X"2B",
X"23",
X"E7",
X"CB",
X"D5",
X"0E",
X"32",
X"25",
X"F7",
X"CB",
X"D5",
X"01",
X"2E",
X"1F",
X"00",
X"CA",
X"DD",
X"FE",
X"31",
X"1B",
X"03",
X"C3",
X"E0",
X"F7",
X"3A",
X"1E",
X"09",
X"BF",
X"DC",
X"EB",
X"3D",
X"1F",
X"15",
X"C3",
X"DC",
X"E2",
X"38",
X"1A",
X"1B",
X"C7",
X"E0",
X"E4",
X"38",
X"18",
X"1C",
X"C4",
X"DD",
X"E1",
X"38",
X"20",
X"21",
X"C7",
X"D9",
X"D8",
X"31",
X"25",
X"25",
X"D2",
X"D8",
X"D5",
X"29",
X"23",
X"24",
X"DA",
X"D5",
X"D9",
X"24",
X"26",
X"24",
X"DF",
X"CE",
X"D8",
X"1B",
X"2D",
X"28",
X"E8",
X"CC",
X"D6",
X"0E",
X"30",
X"27",
X"F4",
X"CF",
X"D8",
X"06",
X"31",
X"1F",
X"FB",
X"CB",
X"DB",
X"02",
X"35",
X"20",
X"00",
X"C3",
X"DA",
X"FB",
X"38",
X"24",
X"0A",
X"C2",
X"D8",
X"EF",
X"37",
X"24",
X"13",
X"C8",
X"DC",
X"E7",
X"34",
X"1F",
X"17",
X"CB",
X"DD",
X"E6",
X"36",
X"1F",
X"1B",
X"CA",
X"D8",
X"E1",
X"33",
X"24",
X"23",
X"CE",
X"D6",
X"D9",
X"2A",
X"25",
X"26",
X"D6",
X"D8",
X"D9",
X"25",
X"26",
X"23",
X"DB",
X"D5",
X"D9",
X"23",
X"2A",
X"25",
X"E1",
X"CF",
X"D6",
X"1B",
X"2E",
X"29",
X"EC",
X"CE",
X"D5",
X"0F",
X"2D",
X"27",
X"F3",
X"CF",
X"DA",
X"08",
X"2F",
X"23",
X"F8",
X"CC",
X"D9",
X"04",
X"34",
X"24",
X"00",
X"C8",
X"D7",
X"FC",
X"35",
X"25",
X"0A",
X"CA",
X"D9",
X"F3",
X"31",
X"21",
X"0E",
X"CC",
X"DD",
X"EF",
X"33",
X"21",
X"11",
X"CB",
X"DB",
X"E9",
X"33",
X"24",
X"18",
X"CD",
X"D8",
X"E2",
X"2F",
X"24",
X"20",
X"D3",
X"D8",
X"DF",
X"29",
X"22",
X"22",
X"D7",
X"DA",
X"DE",
X"26",
X"24",
X"22",
X"DA",
X"D7",
X"D9",
X"22",
X"28",
X"25",
X"E0",
X"D5",
X"D6",
X"1A",
X"28",
X"27",
X"E9",
X"D4",
X"D7",
X"13",
X"27",
X"25",
X"EF",
X"D2",
X"D9",
X"0E",
X"2B",
X"25",
X"F3",
X"CF",
X"D8",
X"06",
X"2F",
X"26",
X"FD",
X"CE",
X"D6",
X"FF",
X"30",
X"25",
X"04",
X"CF",
X"D9",
X"F8",
X"2E",
X"21",
X"0B",
X"CD",
X"DC",
X"F3",
X"30",
X"21",
X"0F",
X"CB",
X"DC",
X"EB",
X"31",
X"22",
X"17",
X"CF",
X"DB",
X"E2",
X"2E",
X"1F",
X"1E",
X"D3",
X"DD",
X"DF",
X"2B",
X"1D",
X"20",
X"D4",
X"DD",
X"DD",
X"29",
X"1F",
X"23",
X"D5",
X"DB",
X"D8",
X"25",
X"22",
X"28",
X"DC",
X"DA",
X"D4",
X"1E",
X"21",
X"29",
X"E5",
X"DB",
X"D5",
X"18",
X"21",
X"27",
X"E9",
X"D9",
X"D7",
X"14",
X"25",
X"26",
X"EE",
X"D4",
X"D6",
X"0B",
X"2A",
X"27",
X"F8",
X"D2",
X"D8",
X"05",
X"2A",
X"25",
X"01",
X"DA",
X"DF",
X"FF",
X"29",
X"1F",
X"07",
X"D6",
X"E2",
X"F9",
X"2C",
X"1D",
X"0D",
X"D3",
X"E1",
X"F0",
X"2E",
X"1D",
X"15",
X"D2",
X"E2",
X"E6",
X"2B",
X"19",
X"1B",
X"D4",
X"E4",
X"E1",
X"29",
X"16",
X"1F",
X"D5",
X"E5",
X"DD",
X"29",
X"17",
X"22",
X"D5",
X"E3",
X"D8",
X"26",
X"18",
X"25",
X"DA",
X"E2",
X"D5",
X"20",
X"18",
X"28",
X"E0",
X"E2",
X"D4",
X"1A",
X"19",
X"27",
X"E6",
X"E0",
X"D5",
X"14",
X"1C",
X"26",
X"EB",
X"DC",
X"D6",
X"0D",
X"1F",
X"24",
X"F3",
X"D9",
X"D6",
X"05",
X"22",
X"23",
X"FD",
X"D8",
X"D9",
X"FE",
X"24",
X"1F",
X"03",
X"D6",
X"DD",
X"F7",
X"28",
X"1C",
X"0A",
X"D2",
X"DF",
X"F0",
X"2A",
X"1B",
X"12",
X"D1",
X"E0",
X"E8",
X"2B",
X"19",
X"19",
X"D2",
X"E2",
X"E2",
X"2A",
X"17",
X"1E",
X"D3",
X"E4",
X"DE",
X"2A",
X"18",
X"22",
X"D5",
X"E3",
X"D9",
X"27",
X"19",
X"25",
X"DA",
X"E3",
X"D6",
X"21",
X"19",
X"27",
X"DF",
X"E2",
X"D6",
X"1C",
X"1A",
X"26",
X"E5",
X"E0",
X"D8",
X"17",
X"1E",
X"26",
X"EC",
X"DC",
X"D7",
X"10",
X"21",
X"26",
X"F5",
X"DB",
X"D9",
X"06",
X"23",
X"23",
X"FD",
X"D9",
X"DC",
X"00",
X"26",
X"20",
X"01",
X"D5",
X"DE",
X"FB",
X"29",
X"1E",
X"09",
X"D3",
X"DE",
X"F2",
X"2B",
X"1E",
X"12",
X"D4",
X"E0",
X"EB",
X"2A",
X"1B",
X"18",
X"D5",
X"E2",
X"E7",
X"2A",
X"1A",
X"1C",
X"D5",
X"E2",
X"E2",
X"29",
X"1C",
X"21",
X"D8",
X"E1",
X"DD",
X"26",
X"1C",
X"24",
X"DD",
X"E1",
X"DB",
X"20",
X"1C",
X"26",
X"E2",
X"E0",
X"DB",
X"1C",
X"1F",
X"25",
X"E7",
X"DE",
X"D9",
X"17",
X"22",
X"26",
X"EE",
X"DB",
X"D8",
X"0F",
X"24",
X"27",
X"F6",
X"D9",
X"DA",
X"08",
X"25",
X"25",
X"FC",
X"D8",
X"DB",
X"01",
X"27",
X"23",
X"01",
X"D6",
X"DC",
X"FC",
X"2A",
X"22",
X"08",
X"D4",
X"DD",
X"F5",
X"2B",
X"20",
X"0F",
X"D5",
X"DE",
X"EF",
X"2A",
X"1F",
X"15",
X"D5",
X"E0",
X"E9",
X"29",
X"1D",
X"19",
X"D6",
X"E0",
X"E5",
X"29",
X"1E",
X"1E",
X"D8",
X"DF",
X"E1",
X"26",
X"1E",
X"23",
X"DC",
X"DF",
X"DD",
X"22",
X"1E",
X"24",
X"E0",
X"DF",
X"DB",
X"1E",
X"1F",
X"25",
X"E4",
X"DE",
X"DA",
X"19",
X"21",
X"27",
X"EA",
X"DB",
X"D8",
X"14",
X"23",
X"28",
X"F1",
X"DB",
X"D8",
X"0D",
X"23",
X"27",
X"F8",
X"D9",
X"D9",
X"07",
X"25",
X"25",
X"FE",
X"D8",
X"DA",
X"00",
X"28",
X"24",
X"02",
X"D6",
X"DA",
X"FB",
X"29",
X"24",
X"0A",
X"D6",
X"DB",
X"F4",
X"29",
X"22",
X"10",
X"D5",
X"DD",
X"EE",
X"2A",
X"20",
X"16",
X"D5",
X"DE",
X"E9",
X"2A",
X"20",
X"1B",
X"D6",
X"DE",
X"E3",
X"29",
X"1F",
X"20",
X"D9",
X"DF",
X"DE",
X"26",
X"1E",
X"24",
X"DB",
X"DF",
X"DB",
X"23",
X"1E",
X"27",
X"DE",
X"DF",
X"D8",
X"1F",
X"1F",
X"29",
X"E3",
X"DE",
X"D6",
X"1A",
X"20",
X"2A",
X"E9",
X"DD",
X"D5",
X"15",
X"21",
X"2A",
X"EE",
X"DC",
X"D4",
X"0E",
X"22",
X"29",
X"F5",
X"DB",
X"D5",
X"08",
X"24",
X"28",
X"FC",
X"D9",
X"D6",
X"01",
X"26",
X"27",
X"01",
X"D6",
X"D7",
X"FB",
X"28",
X"26",
X"08",
X"D5",
X"D9",
X"F4",
X"29",
X"24",
X"0F",
X"D4",
X"DB",
X"ED",
X"2B",
X"22",
X"15",
X"D4",
X"DD",
X"E7",
X"2B",
X"20",
X"1C",
X"D4",
X"DE",
X"E1",
X"2A",
X"1E",
X"21",
X"D6",
X"DF",
X"DB",
X"28",
X"1E",
X"26",
X"D8",
X"DF",
X"D7",
X"25",
X"1D",
X"28",
X"DB",
X"DF",
X"D4",
X"21",
X"1E",
X"2A",
X"E0",
X"DD",
X"D3",
X"1B",
X"20",
X"2C",
X"E6",
X"DC",
X"D2",
X"15",
X"22",
X"2B",
X"ED",
X"DA",
X"D3",
X"0F",
X"24",
X"2A",
X"F4",
X"D7",
X"D4",
X"07",
X"27",
X"28",
X"FC",
X"D5",
X"D6",
X"00",
X"29",
X"25",
X"03",
X"D9",
X"DF",
X"FD",
X"2A",
X"22",
X"09",
X"D6",
X"DF",
X"F5",
X"2B",
X"20",
X"10",
X"D5",
X"E0",
X"EE",
X"2B",
X"1D",
X"16",
X"D4",
X"E2",
X"E8",
X"2B",
X"1B",
X"1B",
X"D5",
X"E2",
X"E1",
X"29",
X"1A",
X"1F",
X"D5",
X"E2",
X"DD",
X"27",
X"1A",
X"22",
X"D8",
X"E1",
X"D9",
X"23",
X"1A",
X"24",
X"DC",
X"DF",
X"D8",
X"1E",
X"1C",
X"24",
X"E1",
X"DD",
X"D7",
X"19",
X"1E",
X"24",
X"E7",
X"DA",
X"D7",
X"12",
X"21",
X"23",
X"EE",
X"D7",
X"D9",
X"0A",
X"24",
X"21",
X"F5",
X"D5",
X"DA",
X"03",
X"27",
X"1F",
X"FD",
X"D2",
X"DC",
X"FE",
X"2A",
X"1D",
X"03",
X"D0",
X"DD",
X"F6",
X"2C",
X"1C",
X"0A",
X"CE",
X"DF",
X"EF",
X"2E",
X"1A",
X"0F",
X"CE",
X"E0",
X"E9",
X"2E",
X"19",
X"15",
X"CE",
X"E1",
X"E5",
X"2D",
X"1A",
X"19",
X"D0",
X"E0",
X"E1",
X"2B",
X"1B",
X"1D",
X"D4",
X"DF",
X"DF",
X"27",
X"1D",
X"1F",
X"D8",
X"DD",
X"DD",
X"22",
X"1E",
X"1F",
X"DD",
X"DB",
X"DC",
X"1D",
X"22",
X"20",
X"E3",
X"D8",
X"DC",
X"16",
X"25",
X"20",
X"EA",
X"D5",
X"DD",
X"10",
X"28",
X"1E",
X"F2",
X"D2",
X"DE",
X"09",
X"2B",
X"1D",
X"F9",
X"D0",
X"DF",
X"02",
X"2E",
X"1C",
X"00",
X"CD",
X"E0",
X"FD",
X"30",
X"1B",
X"04",
X"CC",
X"E1",
X"F6",
X"30",
X"1B",
X"0B",
X"CC",
X"E1",
X"F1",
X"31",
X"1A",
X"10",
X"CC",
X"E1",
X"EC",
X"31",
X"1B",
X"15",
X"CE",
X"E0",
X"E8",
X"2F",
X"1C",
X"18",
X"D0",
X"DF",
X"E4",
X"2B",
X"1E",
X"1B",
X"D4",
X"DE",
X"E2",
X"28",
X"20",
X"1D",
X"D9",
X"DC",
X"E1",
X"23",
X"22",
X"1E",
X"DF",
X"D8",
X"E0",
X"1D",
X"25",
X"1F",
X"E5",
X"D6",
X"DF",
X"17",
X"28",
X"1F",
X"EB",
X"D4",
X"DE",
X"11",
X"2A",
X"1E",
X"F2",
X"D1",
X"DF",
X"0A",
X"2C",
X"1E",
X"F8",
X"CF",
X"DF",
X"03",
X"2E",
X"1E",
X"00",
X"CE",
X"DF",
X"FF",
X"30",
X"1D",
X"04",
X"CE",
X"E0",
X"F8",
X"30",
X"1D",
X"0A",
X"CD",
X"DF",
X"F2",
X"31",
X"1D",
X"10",
X"CE",
X"DF",
X"ED",
X"2F",
X"1D",
X"15",
X"CF",
X"DE",
X"E9",
X"2E",
X"1E",
X"19",
X"D2",
X"DD",
X"E5",
X"2B",
X"1F",
X"1C",
X"D5",
X"DC",
X"E1",
X"28",
X"20",
X"1E",
X"DA",
X"DB",
X"DF",
X"23",
X"23",
X"20",
X"DE",
X"D9",
X"DD",
X"1F",
X"24",
X"22",
X"E4",
X"D7",
X"DC",
X"19",
X"26",
X"22",
X"EA",
X"D5",
X"DB",
X"13",
X"29",
X"22",
X"F1",
X"D3",
X"DB",
X"0C",
X"2B",
X"21",
X"F7",
X"D1",
X"DC",
X"04",
X"2C",
X"21",
X"FE",
X"CF",
X"DC",
X"FF",
X"2E",
X"20",
X"03",
X"CE",
X"DD",
X"F9",
X"2F",
X"1F",
X"0A",
X"CE",
X"DE",
X"F2",
X"30",
X"1F",
X"10",
X"CE",
X"DE",
X"ED",
X"2F",
X"1E",
X"15",
X"D0",
X"DE",
X"E7",
X"2E",
X"1E",
X"19",
X"D2",
X"DE",
X"E3",
X"2B",
X"1F",
X"1D",
X"D5",
X"DD",
X"DF",
X"28",
X"20",
X"20",
X"D9",
X"DB",
X"DD",
X"24",
X"21",
X"22",
X"DF",
X"DA",
X"DC",
X"1E",
X"23",
X"22",
X"E4",
X"D8",
X"DB",
X"18",
X"26",
X"22",
X"EB",
X"D5",
X"DB",
X"10",
X"28",
X"22",
X"F2",
X"D3",
X"DB",
X"09",
X"2A",
X"21",
X"F9",
X"D0",
X"DC",
X"02",
X"2D",
X"20",
X"00",
X"CF",
X"DD",
X"FD",
X"2F",
X"1E",
X"06",
X"CE",
X"DE",
X"F5",
X"30",
X"1D",
X"0D",
X"CD",
X"DF",
X"EF",
X"30",
X"1C",
X"13",
X"CE",
X"E0",
X"E9",
X"2F",
X"1C",
X"18",
X"CF",
X"E0",
X"E4",
X"2D",
X"1C",
X"1C",
X"D3",
X"DE",
X"E0",
X"29",
X"1E",
X"1F",
X"D7",
X"DD",
X"DD",
X"25",
X"1F",
X"20",
X"DB",
X"DB",
X"DC",
X"20",
X"22",
X"21",
X"E1",
X"D8",
X"DC",
X"19",
X"25",
X"21",
X"E9",
X"D5",
X"DC",
X"11",
X"28",
X"21",
X"F1",
X"D2",
X"DC",
X"0A",
X"2B",
X"1F",
X"F9",
X"CF",
X"DE",
X"02",
X"2E",
X"1D",
X"00",
X"CD",
X"DF",
X"FC",
X"30",
X"1C",
X"07",
X"D2",
X"E8",
X"F9",
X"31",
X"19",
X"0D",
X"D1",
X"E7",
X"F3",
X"30",
X"18",
X"11",
X"D0",
X"E7",
X"ED",
X"2F",
X"17",
X"16",
X"D2",
X"E6",
X"E8",
X"2C",
X"17",
X"19",
X"D3",
X"E4",
X"E4",
X"29",
X"18",
X"1A",
X"D7",
X"E3",
X"E1",
X"23",
X"19",
X"1C",
X"DC",
X"E0",
X"DF",
X"1E",
X"1C",
X"1D",
X"E1",
X"DC",
X"DF",
X"18",
X"1F",
X"1C",
X"E8",
X"D9",
X"DF",
X"11",
X"22",
X"1B",
X"EE",
X"D6",
X"DF",
X"09",
X"25",
X"1A",
X"F6",
X"D3",
X"E1",
X"02",
X"28",
X"18",
X"FC",
X"D0",
X"E2",
X"FC",
X"2A",
X"16",
X"02",
X"CF",
X"E3",
X"F6",
X"2C",
X"16",
X"08",
X"CE",
X"E4",
X"F0",
X"2C",
X"15",
X"0E",
X"CF",
X"E4",
X"EB",
X"2C",
X"15",
X"13",
X"D0",
X"E4",
X"E7",
X"2A",
X"16",
X"17",
X"D2",
X"E3",
X"E3",
X"27",
X"17",
X"1A",
X"D6",
X"E2",
X"E0",
X"24",
X"19",
X"1C",
X"DB",
X"E0",
X"DF",
X"1F",
X"1B",
X"1D",
X"E1",
X"DE",
X"DE",
X"19",
X"1E",
X"1E",
X"E6",
X"DB",
X"DE",
X"13",
X"21",
X"1D",
X"ED",
X"D9",
X"DE",
X"0D",
X"23",
X"1C",
X"F4",
X"D7",
X"E0",
X"06",
X"26",
X"1C",
X"FB",
X"D5",
X"E0",
X"00",
X"28",
X"1B",
X"00",
X"D4",
X"E1",
X"FB",
X"29",
X"1A",
X"06",
X"D4",
X"E2",
X"F5",
X"29",
X"1A",
X"0C",
X"D3",
X"E2",
X"EF",
X"29",
X"19",
X"11",
X"D4",
X"E2",
X"EA",
X"28",
X"1A",
X"16",
X"D6",
X"E2",
X"E6",
X"26",
X"1A",
X"19",
X"D9",
X"E1",
X"E3",
X"24",
X"1B",
X"1C",
X"DD",
X"E0",
X"E0",
X"20",
X"1D",
X"1E",
X"E1",
X"E0",
X"DE",
X"1B",
X"1E",
X"21",
X"E6",
X"DE",
X"DD",
X"16",
X"20",
X"21",
X"EC",
X"DC",
X"DC",
X"10",
X"21",
X"22",
X"F2",
X"DB",
X"DC",
X"0A",
X"23",
X"21",
X"F8",
X"DA",
X"DC",
X"04",
X"24",
X"21",
X"FE",
X"D8",
X"DC",
X"FF",
X"25",
X"20",
X"03",
X"D8",
X"DD",
X"F9",
X"26",
X"1F",
X"09",
X"D8",
X"DE",
X"F3",
X"27",
X"1E",
X"0F",
X"D8",
X"DE",
X"ED",
X"26",
X"1D",
X"14",
X"D9",
X"DF",
X"E8",
X"25",
X"1D",
X"19",
X"DB",
X"E0",
X"E4",
X"23",
X"1C",
X"1D",
X"DD",
X"E0",
X"E0",
X"20",
X"1C",
X"20",
X"E1",
X"E0",
X"DD",
X"1C",
X"1D",
X"22",
X"E5",
X"DF",
X"DB",
X"18",
X"1E",
X"24",
X"EA",
X"DE",
X"D9",
X"13",
X"1F",
X"24",
X"EF",
X"DD",
X"D9",
X"0D",
X"21",
X"24",
X"F5",
X"DC",
X"DA",
X"07",
X"22",
X"24",
X"FC",
X"DB",
X"DA",
X"00",
X"23",
X"23",
X"01",
X"DA",
X"DB",
X"FC",
X"24",
X"21",
X"07",
X"D9",
X"DC",
X"F5",
X"26",
X"1F",
X"0E",
X"D8",
X"DE",
X"EE",
X"26",
X"1E",
X"14",
X"D8",
X"DF",
X"E8",
X"25",
X"1C",
X"1A",
X"D9",
X"E1",
X"E3",
X"24",
X"1C",
X"1E",
X"DB",
X"E1",
X"DE",
X"22",
X"1B",
X"22",
X"DE",
X"E1",
X"DB",
X"1E",
X"1B",
X"25",
X"E2",
X"E0",
X"D8",
X"1A",
X"1D",
X"26",
X"E7",
X"DF",
X"D7",
X"15",
X"1E",
X"27",
X"ED",
X"DE",
X"D7",
X"0F",
X"1F",
X"26",
X"F3",
X"DC",
X"D7",
X"08",
X"21",
X"25",
X"FA",
X"DA",
X"D8",
X"01",
X"24",
X"24",
X"00",
X"D8",
X"DA",
X"FB",
X"26",
X"22",
X"07",
X"D6",
X"DC",
X"F4",
X"27",
X"1F",
X"0E",
X"D5",
X"DE",
X"ED",
X"28",
X"1D",
X"15",
X"D5",
X"E0",
X"E7",
X"28",
X"1B",
X"1B",
X"D6",
X"E1",
X"E1",
X"27",
X"1A",
X"20",
X"D8",
X"E2",
X"DD",
X"24",
X"1A",
X"23",
X"DA",
X"E2",
X"D9",
X"21",
X"1A",
X"27",
X"DE",
X"E2",
X"D7",
X"1D",
X"1A",
X"28",
X"E4",
X"E0",
X"D6",
X"18",
X"1D",
X"28",
X"EA",
X"DE",
X"D6",
X"11",
X"1E",
X"27",
X"F0",
X"DC",
X"D6",
X"0A",
X"21",
X"25",
X"F7",
X"D9",
X"D8",
X"03",
X"23",
X"23",
X"FE",
X"D7",
X"DA",
X"FD",
X"26",
X"21",
X"04",
X"D5",
X"DC",
X"F6",
X"27",
X"1F",
X"0C",
X"D4",
X"DE",
X"EF",
X"29",
X"1C",
X"13",
X"D3",
X"E5",
X"EE",
X"28",
X"1B",
X"18",
X"DA",
X"E7",
X"E8",
X"27",
X"19",
X"1C",
X"DA",
X"E7",
X"E3",
X"25",
X"17",
X"1F",
X"DC",
X"E7",
X"DF",
X"21",
X"17",
X"21",
X"DF",
X"E6",
X"DC",
X"1D",
X"18",
X"22",
X"E3",
X"E4",
X"DB",
X"18",
X"19",
X"22",
X"E8",
X"E1",
X"DA",
X"12",
X"1A",
X"22",
X"ED",
X"DF",
X"DA",
X"0C",
X"1C",
X"21",
X"F3",
X"DD",
X"DB",
X"05",
X"1D",
X"1F",
X"FA",
X"DB",
X"DC",
X"00",
X"20",
X"1D",
X"00",
X"DA",
X"DD",
X"FA",
X"21",
X"1C",
X"04",
X"D8",
X"DE",
X"F4",
X"22",
X"1A",
X"09",
X"D7",
X"E0",
X"EF",
X"22",
X"19",
X"0F",
X"D7",
X"E0",
X"EA",
X"22",
X"18",
X"14",
X"DA",
X"E1",
X"E6",
X"21",
X"18",
X"17",
X"DB",
X"E1",
X"E2",
X"1F",
X"19",
X"1B",
X"DD",
X"E1",
X"E0",
X"1C",
X"19",
X"1D",
X"E1",
X"E0",
X"DE",
X"19",
X"1A",
X"1F",
X"E5",
X"DF",
X"DD",
X"15",
X"1C",
X"1F",
X"EA",
X"DF",
X"DC",
X"10",
X"1D",
X"1F",
X"F0",
X"DD",
X"DC",
X"0B",
X"1F",
X"1F",
X"F5",
X"DC",
X"DC",
X"06",
X"20",
X"1F",
X"FA",
X"DB",
X"DD",
X"00",
X"21",
X"1E",
X"00",
X"DA",
X"DE",
X"FD",
X"22",
X"1E",
X"03",
X"D9",
X"DE",
X"F7",
X"23",
X"1D",
X"09",
X"DA",
X"DF",
X"F3",
X"23",
X"1D",
X"0E",
X"DA",
X"DF",
X"EE",
X"23",
X"1C",
X"12",
X"DB",
X"E0",
X"EA",
X"21",
X"1C",
X"15",
X"DD",
X"E0",
X"E7",
X"1F",
X"1C",
X"19",
X"E0",
X"E0",
X"E4",
X"1D",
X"1C",
X"1B",
X"E3",
X"E0",
X"E1",
X"1A",
X"1D",
X"1E",
X"E7",
X"E0",
X"DF",
X"16",
X"1D",
X"1F",
X"EB",
X"DF",
X"DE",
X"12",
X"1F",
X"20",
X"F0",
X"DE",
X"DE",
X"0D",
X"20",
X"20",
X"F5",
X"DD",
X"DE",
X"08",
X"22",
X"1F",
X"FB",
X"DC",
X"DE",
X"02",
X"23",
X"1F",
X"00",
X"DB",
X"DE",
X"FE",
X"24",
X"1E",
X"04",
X"D9",
X"E0",
X"F8",
X"24",
X"1D",
X"09",
X"D9",
X"E0",
X"F3",
X"24",
X"1C",
X"0F",
X"D9",
X"E1",
X"EE",
X"25",
X"1B",
X"13",
X"DA",
X"E2",
X"E9",
X"24",
X"1A",
X"18",
X"DB",
X"E2",
X"E5",
X"23",
X"1A",
X"1B",
X"DD",
X"E3",
X"E2",
X"20",
X"1A",
X"1E",
X"E1",
X"E2",
X"DF",
X"1D",
X"1B",
X"20",
X"E5",
X"E1",
X"DE",
X"19",
X"1C",
X"20",
X"E9",
X"E0",
X"DD",
X"14",
X"1E",
X"21",
X"EF",
X"DE",
X"DD",
X"0E",
X"20",
X"20",
X"F4",
X"DC",
X"DE",
X"08",
X"22",
X"1F",
X"FB",
X"DA",
X"E0",
X"01",
X"25",
X"1D",
X"00",
X"D8",
X"E1",
X"FD",
X"27",
X"1B",
X"06",
X"D7",
X"E2",
X"F6",
X"28",
X"19",
X"0C",
X"D6",
X"E4",
X"F0",
X"29",
X"18",
X"11",
X"D5",
X"E6",
X"EB",
X"29",
X"17",
X"16",
X"D5",
X"E6",
X"E6",
X"28",
X"16",
X"1A",
X"D7",
X"E6",
X"E3",
X"26",
X"17",
X"1C",
X"DA",
X"E6",
X"E1",
X"23",
X"18",
X"1E",
X"DF",
X"E5",
X"DF",
X"1F",
X"19",
X"1F",
X"E3",
X"E3",
X"DE",
X"19",
X"1C",
X"1F",
X"E8",
X"E0",
X"DE",
X"14",
X"1F",
X"1E",
X"EE",
X"DD",
X"E0",
X"0D",
X"21",
X"1D",
X"F5",
X"DA",
X"E1",
X"06",
X"24",
X"1B",
X"FC",
X"D8",
X"E2",
X"00",
X"27",
X"19",
X"01",
X"D5",
X"E4",
X"FB",
X"28",
X"18",
X"07",
X"D4",
X"E6",
X"F5",
X"2A",
X"17",
X"0D",
X"D3",
X"E6",
X"EF",
X"2B",
X"16",
X"12",
X"D4",
X"E7",
X"EB",
X"2A",
X"15",
X"16",
X"D5",
X"E7",
X"E7",
X"29",
X"16",
X"19",
X"D7",
X"E6",
X"E4",
X"25",
X"17",
X"1B",
X"DB",
X"E4",
X"E3",
X"20",
X"19",
X"1C",
X"DF",
X"E3",
X"E1",
X"1C",
X"1B",
X"1D",
X"E5",
X"E0",
X"E1",
X"17",
X"1E",
X"1C",
X"EB",
X"DD",
X"E2",
X"11",
X"21",
X"1B",
X"F0",
X"DA",
X"E2",
X"0A",
X"23",
X"1A",
X"F7",
X"D7",
X"E4",
X"03",
X"26",
X"18",
X"FE",
X"D5",
X"E5",
X"FF",
X"27",
X"17",
X"02",
X"D4",
X"E5",
X"F9",
X"29",
X"16",
X"07",
X"D4",
X"E6",
X"F4",
X"29",
X"16",
X"0D",
X"DB",
X"ED",
X"F6",
X"28",
X"15",
X"0F",
X"DB",
X"EC",
X"F1",
X"25",
X"15",
X"11",
X"DC",
X"EA",
X"EE",
X"23",
X"15",
X"13",
X"DE",
X"E8",
X"EC",
X"1F",
X"16",
X"14",
X"E1",
X"E6",
X"EA",
X"1B",
X"18",
X"14",
X"E5",
X"E4",
X"E8",
X"16",
X"1A",
X"14",
X"E9",
X"E1",
X"E8",
X"10",
X"1B",
X"13",
X"ED",
X"DE",
X"E8",
X"0C",
X"1D",
X"13",
X"F2",
X"DC",
X"E8",
X"06",
X"1F",
X"12",
X"F8",
X"DA",
X"E7",
X"01",
X"20",
X"12",
X"FC",
X"D9",
X"E8",
X"FE",
X"21",
X"12",
X"00",
X"D8",
X"E8",
X"FA",
X"22",
X"12",
X"03",
X"D8",
X"E8",
X"F6",
X"22",
X"12",
X"08",
X"D9",
X"E7",
X"F2",
X"21",
X"13",
X"0B",
X"DA",
X"E6",
X"EF",
X"20",
X"13",
X"0D",
X"DC",
X"E6",
X"EC",
X"1E",
X"15",
X"10",
X"DF",
X"E4",
X"EB",
X"1B",
X"17",
X"12",
X"E2",
X"E3",
X"E9",
X"18",
X"18",
X"13",
X"E6",
X"E1",
X"E8",
X"14",
X"1A",
X"14",
X"EA",
X"E0",
X"E8",
X"10",
X"1C",
X"14",
X"EF",
X"DE",
X"E8",
X"0B",
X"1E",
X"14",
X"F4",
X"DD",
X"E8",
X"06",
X"20",
X"15",
X"F9",
X"DC",
X"E8",
X"02",
X"21",
X"14",
X"FF",
X"DB",
X"E8",
X"FF",
X"22",
X"14",
X"01",
X"DA",
X"E8",
X"FA",
X"23",
X"13",
X"06",
X"DA",
X"E9",
X"F5",
X"23",
X"13",
X"0A",
X"DA",
X"E9",
X"F1",
X"23",
X"14",
X"0E",
X"DB",
X"E8",
X"ED",
X"21",
X"14",
X"12",
X"DD",
X"E7",
X"EA",
X"1F",
X"15",
X"15",
X"E0",
X"E7",
X"E8",
X"1D",
X"16",
X"17",
X"E3",
X"E5",
X"E6",
X"1A",
X"18",
X"19",
X"E8",
X"E4",
X"E5",
X"15",
X"1A",
X"19",
X"EC",
X"E2",
X"E5",
X"10",
X"1C",
X"19",
X"F2",
X"E0",
X"E5",
X"0B",
X"1E",
X"18",
X"F7",
X"DE",
X"E6",
X"05",
X"20",
X"18",
X"FD",
X"DD",
X"E6",
X"00",
X"22",
X"17",
X"00",
X"DB",
X"E7",
X"FB",
X"23",
X"15",
X"06",
X"D9",
X"E8",
X"F5",
X"24",
X"14",
X"0B",
X"D9",
X"E9",
X"F0",
X"24",
X"14",
X"10",
X"DA",
X"EA",
X"EC",
X"24",
X"13",
X"15",
X"DB",
X"EA",
X"E8",
X"23",
X"14",
X"18",
X"DD",
X"E9",
X"E5",
X"20",
X"15",
X"1A",
X"E0",
X"E8",
X"E4",
X"1D",
X"16",
X"1C",
X"E4",
X"E7",
X"E3",
X"18",
X"17",
X"1C",
X"E9",
X"E5",
X"E1",
X"13",
X"1A",
X"1C",
X"EF",
X"E3",
X"E2",
X"0D",
X"1C",
X"1B",
X"F5",
X"E0",
X"E3",
X"07",
X"1F",
X"1A",
X"FB",
X"DE",
X"E4",
X"01",
X"21",
X"18",
X"00",
X"DB",
X"E6",
X"FC",
X"23",
X"17",
X"06",
X"DA",
X"E7",
X"F6",
X"25",
X"15",
X"0B",
X"D9",
X"E8",
X"F0",
X"25",
X"14",
X"11",
X"D9",
X"E8",
X"EC",
X"25",
X"14",
X"15",
X"DB",
X"E9",
X"E8",
X"23",
X"14",
X"18",
X"DC",
X"E8",
X"E5",
X"21",
X"15",
X"1B",
X"E0",
X"E7",
X"E3",
X"1D",
X"16",
X"1C",
X"E4",
X"E6",
X"E2",
X"19",
X"18",
X"1C",
X"E9",
X"E4",
X"E1",
X"13",
X"1B",
X"1C",
X"EF",
X"E2",
X"E2",
X"0D",
X"1D",
X"1C",
X"F4",
X"DF",
X"E2",
X"08",
X"1F",
X"1A",
X"FB",
X"DD",
X"E3",
X"01",
X"21",
X"19",
X"00",
X"DB",
X"E4",
X"FD",
X"23",
X"18",
X"05",
X"DA",
X"E5",
X"F6",
X"24",
X"17",
X"0B",
X"D9",
X"E6",
X"F1",
X"24",
X"17",
X"0F",
X"DA",
X"E6",
X"ED",
X"23",
X"16",
X"13",
X"DB",
X"E6",
X"E9",
X"22",
X"17",
X"17",
X"DE",
X"E5",
X"E6",
X"1F",
X"17",
X"1A",
X"E1",
X"E5",
X"E3",
X"1C",
X"19",
X"1B",
X"E5",
X"E3",
X"E2",
X"17",
X"1A",
X"1C",
X"E9",
X"E1",
X"E1",
X"12",
X"1C",
X"1C",
X"EF",
X"DE",
X"E1",
X"0C",
X"1E",
X"1B",
X"F5",
X"DD",
X"E2",
X"07",
X"20",
X"1B",
X"FA",
X"DB",
X"E2",
X"01",
X"22",
X"1A",
X"00",
X"DA",
X"E2",
X"FD",
X"23",
X"1A",
X"04",
X"D9",
X"E3",
X"F7",
X"23",
X"19",
X"09",
X"D9",
X"E2",
X"F2",
X"23",
X"19",
X"0E",
X"D9",
X"E2",
X"EE",
X"23",
X"19",
X"12",
X"DB",
X"E2",
X"E9",
X"21",
X"19",
X"16",
X"E5",
X"EB",
X"ED",
X"1E",
X"18",
X"17",
X"E6",
X"E9",
X"EA",
X"1A",
X"18",
X"18",
X"E9",
X"E8",
X"E7",
X"16",
X"17",
X"19",
X"EC",
X"E6",
X"E6",
X"12",
X"17",
X"19",
X"EF",
X"E5",
X"E4",
X"0D",
X"19",
X"19",
X"F3",
X"E3",
X"E3",
X"08",
X"1B",
X"19",
X"F7",
X"E0",
X"E2",
X"03",
X"1B",
X"19",
X"FC",
X"DF",
X"E2",
X"FF",
X"1C",
X"18",
X"00",
X"DD",
X"E3",
X"FA",
X"1C",
X"17",
X"03",
X"DD",
X"E3",
X"F5",
X"1C",
X"16",
X"08",
X"DD",
X"E3",
X"F0",
X"1D",
X"16",
X"0C",
X"DD",
X"E4",
X"EC",
X"1C",
X"15",
X"10",
X"DE",
X"E5",
X"E9",
X"1A",
X"15",
X"14",
X"E1",
X"E4",
X"E5",
X"19",
X"15",
X"17",
X"E3",
X"E4",
X"E3",
X"17",
X"15",
X"19",
X"E6",
X"E5",
X"E1",
X"14",
X"16",
X"1A",
X"E9",
X"E4",
X"E0",
X"10",
X"17",
X"1C",
X"EE",
X"E4",
X"DF",
X"0C",
X"18",
X"1D",
X"F2",
X"E4",
X"DF",
X"08",
X"19",
X"1D",
X"F8",
X"E2",
X"E0",
X"03",
X"1A",
X"1C",
X"FD",
X"E1",
X"E0",
X"00",
X"1B",
X"1C",
X"00",
X"E0",
X"E1",
X"FA",
X"1C",
X"1A",
X"05",
X"E0",
X"E3",
X"F6",
X"1D",
X"19",
X"0A",
X"DF",
X"E4",
X"F1",
X"1D",
X"18",
X"0F",
X"DF",
X"E5",
X"EC",
X"1D",
X"17",
X"13",
X"E0",
X"E6",
X"E8",
X"1C",
X"16",
X"17",
X"E1",
X"E7",
X"E4",
X"1B",
X"15",
X"1A",
X"E3",
X"E7",
X"E2",
X"19",
X"16",
X"1D",
X"E6",
X"E7",
X"E0",
X"15",
X"16",
X"1E",
X"EA",
X"E7",
X"DF",
X"12",
X"17",
X"1F",
X"EF",
X"E6",
X"DF",
X"0E",
X"18",
X"1F",
X"F3",
X"E4",
X"DF",
X"08",
X"1A",
X"1F",
X"F9",
X"E3",
X"E0",
X"03",
X"1B",
X"1E",
X"FF",
X"E1",
X"E1",
X"FF",
X"1D",
X"1C",
X"03",
X"E0",
X"E3",
X"F9",
X"1E",
X"1A",
X"08",
X"DF",
X"E4",
X"F4",
X"1F",
X"19",
X"0D",
X"DF",
X"E5",
X"EE",
X"1F",
X"17",
X"12",
X"DF",
X"E6",
X"EA"  );
--//--------------------------------------
  begin

    if (RESET_N='0') then
      Q <= sqr_table(0);
    elsif(rising_edge(CLK)) then
      if (ENA='1') then
          Q <= sqr_table(to_integer(unsigned(ADDR)));
      end if;
    end if;
  end process;
end arch;