
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.std_logic_unsigned.all;
use ieee.numeric_std.all;
-- Saar Eliad 2017 

entity background is
port 	(
		--////////////////////	Clock Input	 	////////////////////	
	   CLK  : in std_logic;
		RESETn	: in std_logic;
		oCoord_X 		: in integer;
		oCoord_Y 		: in integer;
		mVGA_RGB	      : out std_logic_vector(7 downto 0) --	,   						//	VGA Red[9:0]

	);
end entity;

architecture arch_background of background is 


signal mVGA_R	: std_logic_vector(2 downto 0); --	,	 						//	VGA Red[9:0]
signal mVGA_G	: std_logic_vector(2 downto 0); --	,	 						//	VGA Green[9:0]
signal mVGA_B	:  std_logic_vector(1 downto 0); --	,  						//	VGA Blue[9:0]
	
begin

mVGA_RGB <=  mVGA_R & mVGA_G &  mVGA_B ;

mVGA_R <= "111" when (oCoord_y >= 256 and oCoord_X > 156) else
			 "110" ;	
mVGA_G <= "111" when (oCoord_X <  356 and oCoord_Y < 100) else
 		    "110" ;	
mVGA_B <= "10" when (oCoord_X <  300 and oCoord_Y < 200) else
			 "00";	 
		
end architecture;		