--------------------------------------
-- SinTable.vhd
-- Written by Saar Eliad and Itamar Raviv.
-- All rights reserved, Copyright 2017
--------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity JumpSoundTable is
port(
  CLK     : in std_logic;
  RESET_N : in std_logic;
  ENA     : in std_logic;
  ADDR    : in std_logic_vector(11 downto 0);
  Q       : out std_logic_vector(7 downto 0)
);
end JumpSoundTable;

architecture arch of JumpSoundTable is

type table_type is array(0 to 4095) of std_logic_vector(7 downto 0);
signal sqr_table : table_type;

begin

  JumpSoundTable_proc: process(RESET_N, CLK)
    constant sqr_table : table_type := (
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"01",
X"00",
X"00",
X"FF",
X"00",
X"FE",
X"01",
X"FF",
X"01",
X"FD",
X"00",
X"FF",
X"00",
X"FF",
X"01",
X"FF",
X"00",
X"00",
X"00",
X"FD",
X"01",
X"FE",
X"01",
X"FF",
X"01",
X"FD",
X"00",
X"FC",
X"00",
X"FC",
X"02",
X"FB",
X"04",
X"FB",
X"08",
X"F5",
X"3F",
X"7D",
X"73",
X"73",
X"73",
X"6D",
X"74",
X"69",
X"7A",
X"3D",
X"EE",
X"FC",
X"F7",
X"FA",
X"F9",
X"F8",
X"FC",
X"F3",
X"18",
X"76",
X"68",
X"6D",
X"66",
X"68",
X"66",
X"66",
X"6A",
X"51",
X"EB",
X"F4",
X"EE",
X"F4",
X"EF",
X"F2",
X"F1",
X"F2",
X"FA",
X"64",
X"64",
X"66",
X"60",
X"64",
X"62",
X"64",
X"5E",
X"5D",
X"F5",
X"EA",
X"EA",
X"EC",
X"E8",
X"ED",
X"E7",
X"F1",
X"E6",
X"4A",
X"63",
X"5B",
X"5C",
X"5F",
X"5B",
X"5E",
X"54",
X"62",
X"07",
X"DD",
X"E7",
X"E2",
X"E2",
X"E5",
X"E2",
X"E9",
X"DA",
X"27",
X"63",
X"54",
X"5A",
X"56",
X"55",
X"57",
X"52",
X"5E",
X"1E",
X"D3",
X"E4",
X"DB",
X"E0",
X"DD",
X"DF",
X"E2",
X"D6",
X"04",
X"5E",
X"4F",
X"53",
X"46",
X"4D",
X"48",
X"48",
X"4D",
X"30",
X"D3",
X"E0",
X"D7",
X"E0",
X"D7",
X"DE",
X"DB",
X"DB",
X"E8",
X"4C",
X"44",
X"4B",
X"43",
X"4A",
X"44",
X"47",
X"41",
X"41",
X"DC",
X"D8",
X"D6",
X"DB",
X"D5",
X"DB",
X"D5",
X"DC",
X"D3",
X"35",
X"46",
X"45",
X"43",
X"46",
X"40",
X"46",
X"3D",
X"4A",
X"EF",
X"CE",
X"D3",
X"D3",
X"D3",
X"D5",
X"D0",
X"D9",
X"C9",
X"17",
X"4B",
X"40",
X"43",
X"3E",
X"3F",
X"41",
X"38",
X"47",
X"06",
X"C4",
X"D3",
X"CB",
X"D1",
X"D0",
X"CF",
X"D5",
X"C8",
X"F9",
X"4A",
X"3A",
X"42",
X"3B",
X"3D",
X"3C",
X"3A",
X"3F",
X"1D",
X"C2",
X"D1",
X"C8",
X"D1",
X"CB",
X"CE",
X"CC",
X"CD",
X"E0",
X"41",
X"37",
X"3F",
X"37",
X"3D",
X"36",
X"3A",
X"37",
X"31",
X"CB",
X"CB",
X"C8",
X"CC",
X"C7",
X"CF",
X"C8",
X"CE",
X"CB",
X"29",
X"33",
X"33",
X"2F",
X"32",
X"2C",
X"32",
X"29",
X"34",
X"DC",
X"C4",
X"C8",
X"CA",
X"C8",
X"CC",
X"C7",
X"CF",
X"C2",
X"12",
X"37",
X"2D",
X"31",
X"2F",
X"2D",
X"31",
X"29",
X"36",
X"F5",
X"BC",
X"CB",
X"C4",
X"C9",
X"C6",
X"C6",
X"CA",
X"C1",
X"F1",
X"3B",
X"2A",
X"33",
X"2C",
X"31",
X"2D",
X"2D",
X"30",
X"13",
X"BC",
X"CA",
X"BF",
X"C9",
X"C4",
X"CB",
X"C6",
X"C7",
X"D0",
X"30",
X"2B",
X"33",
X"29",
X"31",
X"27",
X"2C",
X"27",
X"2C",
X"CB",
X"C5",
X"BF",
X"C6",
X"C0",
X"CB",
X"C1",
X"CB",
X"BE",
X"17",
X"2F",
X"2E",
X"2C",
X"2F",
X"25",
X"2E",
X"24",
X"34",
X"EA",
X"BD",
X"C6",
X"C2",
X"C1",
X"C6",
X"C0",
X"CA",
X"BB",
X"F3",
X"32",
X"20",
X"25",
X"24",
X"24",
X"22",
X"1E",
X"27",
X"05",
X"BC",
X"CA",
X"BF",
X"C4",
X"C0",
X"C4",
X"C1",
X"BD",
X"D1",
X"27",
X"1E",
X"27",
X"22",
X"26",
X"1F",
X"22",
X"1F",
X"1E",
X"C7",
X"C4",
X"C1",
X"C5",
X"BE",
X"C5",
X"C1",
X"C7",
X"C1",
X"1A",
X"27",
X"25",
X"22",
X"25",
X"1F",
X"2A",
X"21",
X"2D",
X"DF",
X"BF",
X"C3",
X"C3",
X"BF",
X"C6",
X"C2",
X"C7",
X"BC",
X"FD",
X"29",
X"22",
X"25",
X"24",
X"22",
X"26",
X"23",
X"2D",
X"FF",
X"BE",
X"C6",
X"C4",
X"C2",
X"C3",
X"BF",
X"C4",
X"B9",
X"E1",
X"3C",
X"36",
X"36",
X"3C",
X"EC",
X"B9",
X"CC",
X"C2",
X"CA",
X"C5",
X"C6",
X"C2",
X"C6",
X"C3",
X"C5",
X"C3",
X"C7",
X"CC",
X"2D",
X"41",
X"37",
X"43",
X"11",
X"B7",
X"C8",
X"BF",
X"C9",
X"C2",
X"CB",
X"C4",
X"CC",
X"C5",
X"CD",
X"C4",
X"CF",
X"BF",
X"11",
X"46",
X"3A",
X"41",
X"2F",
X"CE",
X"C5",
X"C5",
X"C7",
X"C6",
X"C9",
X"C7",
X"CD",
X"C9",
X"CC",
X"C7",
X"D0",
X"C2",
X"F2",
X"46",
X"3C",
X"3F",
X"42",
X"ED",
X"BF",
X"CF",
X"C4",
X"CD",
X"C7",
X"CF",
X"CA",
X"D0",
X"CB",
X"CE",
X"CB",
X"CF",
X"CC",
X"2E",
X"46",
X"3B",
X"47",
X"24",
X"C5",
X"D2",
X"C9",
X"D0",
X"CB",
X"D2",
X"CC",
X"D4",
X"CC",
X"D3",
X"C8",
X"D7",
X"C5",
X"FB",
X"4B",
X"42",
X"40",
X"47",
X"F2",
X"C5",
X"D4",
X"CA",
X"D2",
X"CC",
X"D1",
X"CE",
X"D3",
X"CD",
X"D0",
X"CE",
X"D5",
X"CF",
X"2F",
X"4F",
X"40",
X"4D",
X"2D",
X"CC",
X"D3",
X"CE",
X"D1",
X"D0",
X"D3",
X"CF",
X"D5",
X"D0",
X"D6",
X"CE",
X"D8",
X"C8",
X"F8",
X"4D",
X"46",
X"44",
X"4B",
X"FB",
X"C5",
X"D8",
X"CC",
X"D5",
X"CF",
X"D6",
X"CF",
X"D6",
X"D2",
X"D7",
X"D1",
X"DA",
X"CF",
X"2D",
X"50",
X"45",
X"4E",
X"33",
X"D2",
X"D4",
X"D1",
X"D6",
X"D2",
X"D7",
X"D2",
X"D7",
X"D2",
X"D8",
X"D1",
X"DA",
X"CC",
X"F6",
X"4E",
X"4A",
X"48",
X"4F",
X"01",
X"C8",
X"DB",
X"CF",
X"D9",
X"D1",
X"DB",
X"D3",
X"D9",
X"D5",
X"DB",
X"D3",
X"DC",
X"CF",
X"2C",
X"53",
X"44",
X"50",
X"39",
X"D5",
X"D5",
X"D4",
X"D8",
X"D5",
X"D9",
X"D5",
X"D8",
X"D5",
X"DB",
X"D3",
X"DC",
X"CF",
X"F5",
X"4E",
X"4C",
X"48",
X"53",
X"07",
X"C9",
X"DD",
X"D3",
X"DB",
X"D4",
X"DC",
X"D4",
X"DA",
X"D4",
X"DB",
X"D4",
X"DF",
X"D0",
X"29",
X"57",
X"49",
X"51",
X"3F",
X"DB",
X"D6",
X"D7",
X"D9",
X"D7",
X"DB",
X"D8",
X"DB",
X"D8",
X"DC",
X"D7",
X"DE",
X"D4",
X"F2",
X"4F",
X"50",
X"4B",
X"55",
X"10",
X"CA",
X"DF",
X"D3",
X"DE",
X"D5",
X"DE",
X"D6",
X"DF",
X"D6",
X"DF",
X"D7",
X"E1",
X"D1",
X"27",
X"5A",
X"4B",
X"52",
X"44",
X"E1",
X"D6",
X"DA",
X"DA",
X"DA",
X"DB",
X"DA",
X"DC",
X"DB",
X"DD",
X"DA",
X"E0",
X"D6",
X"EF",
X"4F",
X"53",
X"4C",
X"56",
X"16",
X"CD",
X"E1",
X"D5",
X"E0",
X"D6",
X"DF",
X"D8",
X"E1",
X"D9",
X"E1",
X"D8",
X"E4",
X"D2",
X"23",
X"5B",
X"4D",
X"53",
X"49",
X"E6",
X"D7",
X"DC",
X"DA",
X"DC",
X"DD",
X"DC",
X"DD",
X"DC",
X"DE",
X"DD",
X"E0",
X"D9",
X"ED",
X"4F",
X"56",
X"4F",
X"5A",
X"1D",
X"CF",
X"E2",
X"D6",
X"E1",
X"D9",
X"E1",
X"D9",
X"E2",
X"D9",
X"E2",
X"D9",
X"E6",
X"D3",
X"20",
X"5C",
X"50",
X"55",
X"4D",
X"EB",
X"D7",
X"DF",
X"DB",
X"DF",
X"DD",
X"DE",
X"DD",
X"DF",
X"DF",
X"DF",
X"E0",
X"DD",
X"EB",
X"4D",
X"56",
X"4E",
X"5A",
X"23",
X"D1",
X"E3",
X"D8",
X"E3",
X"DA",
X"E3",
X"DA",
X"E3",
X"DB",
X"E4",
X"DB",
X"E8",
X"D3",
X"1B",
X"5D",
X"50",
X"55",
X"50",
X"F1",
X"D7",
X"E1",
X"DC",
X"E1",
X"DD",
X"E0",
X"DE",
X"E1",
X"DF",
X"E0",
X"E1",
X"DF",
X"E7",
X"4A",
X"59",
X"50",
X"5B",
X"2A",
X"D3",
X"E4",
X"D9",
X"E2",
X"DA",
X"E3",
X"DB",
X"E3",
X"DC",
X"E5",
X"DB",
X"E8",
X"D4",
X"17",
X"5E",
X"51",
X"55",
X"53",
X"F6",
X"D7",
X"E3",
X"DC",
X"E1",
X"DC",
X"E2",
X"DF",
X"E2",
X"E1",
X"E2",
X"E0",
X"E2",
X"E5",
X"49",
X"5B",
X"50",
X"5C",
X"2F",
X"D6",
X"E5",
X"DB",
X"E3",
X"DB",
X"E3",
X"DE",
X"E4",
X"DE",
X"E6",
X"DB",
X"E8",
X"D6",
X"13",
X"5F",
X"53",
X"56",
X"57",
X"FD",
X"D8",
X"E5",
X"DC",
X"E3",
X"DD",
X"E3",
X"E0",
X"E3",
X"E0",
X"E3",
X"DF",
X"E4",
X"E3",
X"45",
X"5B",
X"50",
X"5C",
X"36",
X"D9",
X"E5",
X"DC",
X"E4",
X"DE",
X"E4",
X"DE",
X"E5",
X"DD",
X"E6",
X"DD",
X"EB",
X"D9",
X"0F",
X"5D",
X"54",
X"54",
X"59",
X"01",
X"D7",
X"E6",
X"DC",
X"E5",
X"DF",
X"E5",
X"DF",
X"E4",
X"E0",
X"E4",
X"E0",
X"E8",
X"E1",
X"42",
X"5C",
X"52",
X"5D",
X"3C",
X"DC",
X"E6",
X"DD",
X"E3",
X"DF",
X"E6",
X"DF",
X"E4",
X"E0",
X"E7",
X"DE",
X"EB",
X"DB",
X"09",
X"5E",
X"55",
X"55",
X"5C",
X"07",
X"D6",
X"E8",
X"D9",
X"E4",
X"E0",
X"E7",
X"E0",
X"E8",
X"E0",
X"E4",
X"E1",
X"EA",
X"DF",
X"3F",
X"5F",
X"51",
X"5D",
X"3E",
X"DB",
X"E4",
X"DE",
X"DF",
X"DF",
X"E6",
X"E0",
X"E8",
X"E4",
X"E6",
X"DE",
X"E9",
X"DA",
X"06",
X"5F",
X"57",
X"55",
X"5B",
X"09",
X"D4",
X"E9",
X"DC",
X"E5",
X"E0",
X"E7",
X"DF",
X"E8",
X"E4",
X"E6",
X"E0",
X"E8",
X"E1",
X"3D",
X"62",
X"54",
X"5F",
X"3F",
X"E0",
X"E1",
X"E0",
X"E1",
X"E0",
X"E3",
X"E2",
X"E4",
X"E3",
X"E7",
X"E1",
X"E8",
X"DE",
X"02",
X"5E",
X"59",
X"53",
X"5C",
X"13",
X"D2",
X"E7",
X"DD",
X"E7",
X"DF",
X"E8",
X"E3",
X"E9",
X"E2",
X"E7",
X"DE",
X"E8",
X"D6",
X"1E",
X"63",
X"56",
X"59",
X"57",
X"00",
X"DA",
X"E8",
X"E0",
X"E8",
X"E0",
X"E9",
X"E2",
X"E9",
X"DE",
X"E4",
X"DE",
X"E7",
X"D8",
X"33",
X"60",
X"53",
X"5A",
X"52",
X"F0",
X"E0",
X"E6",
X"DF",
X"E3",
X"E4",
X"E7",
X"E6",
X"E7",
X"E1",
X"E5",
X"E1",
X"E5",
X"E2",
X"43",
X"5E",
X"53",
X"5E",
X"44",
X"E2",
X"E4",
X"E1",
X"E3",
X"E2",
X"E6",
X"E4",
X"E8",
X"E5",
X"E6",
X"E3",
X"E6",
X"E1",
X"EB",
X"32",
X"38",
X"30",
X"3B",
X"1A",
X"DD",
X"E9",
X"E1",
X"E5",
X"E1",
X"E7",
X"E5",
X"EA",
X"E6",
X"E9",
X"E2",
X"EA",
X"E1",
X"FA",
X"37",
X"37",
X"32",
X"3C",
X"0D",
X"DC",
X"EB",
X"E1",
X"E7",
X"E4",
X"E9",
X"E2",
X"EA",
X"E4",
X"EB",
X"E3",
X"ED",
X"DD",
X"09",
X"3D",
X"36",
X"36",
X"3B",
X"00",
X"DF",
X"EC",
X"E4",
X"E9",
X"E4",
X"E8",
X"E4",
X"EB",
X"E5",
X"EB",
X"E6",
X"F0",
X"E1",
X"1A",
X"3F",
X"35",
X"38",
X"36",
X"F2",
X"E4",
X"EC",
X"E7",
X"EA",
X"E7",
X"E8",
X"E6",
X"E9",
X"E9",
X"EC",
X"E9",
X"EC",
X"E6",
X"27",
X"40",
X"35",
X"3C",
X"2C",
X"E9",
X"E9",
X"E9",
X"EA",
X"EA",
X"EA",
X"E8",
X"EB",
X"EB",
X"EB",
X"EA",
X"EC",
X"E8",
X"F0",
X"33",
X"3E",
X"37",
X"3F",
X"22",
X"E5",
X"ED",
X"E7",
X"EC",
X"E8",
X"EC",
X"E8",
X"ED",
X"E9",
X"EE",
X"E9",
X"EF",
X"E4",
X"FC",
X"3B",
X"3C",
X"39",
X"42",
X"15",
X"E1",
X"EF",
X"E6",
X"EE",
X"E7",
X"EC",
X"E8",
X"F0",
X"EA",
X"F0",
X"E8",
X"F1",
X"E3",
X"0A",
X"41",
X"3C",
X"3A",
X"40",
X"06",
X"E2",
X"EF",
X"E6",
X"ED",
X"E9",
X"EE",
X"E9",
X"F1",
X"EA",
X"EF",
X"E8",
X"F3",
X"E4",
X"19",
X"44",
X"3B",
X"3D",
X"3C",
X"FB",
X"E7",
X"EE",
X"E8",
X"ED",
X"EA",
X"EE",
X"EB",
X"EF",
X"EB",
X"EE",
X"EA",
X"F1",
X"E7",
X"28",
X"41",
X"3A",
X"41",
X"34",
X"F0",
X"EC",
X"EC",
X"ED",
X"EE",
X"ED",
X"ED",
X"ED",
X"EE",
X"EC",
X"ED",
X"EE",
X"ED",
X"F0",
X"35",
X"41",
X"3A",
X"42",
X"29",
X"E9",
X"EF",
X"E9",
X"F0",
X"EC",
X"EF",
X"EB",
X"EE",
X"EB",
X"EF",
X"EB",
X"F2",
X"EA",
X"FD",
X"3F",
X"41",
X"3C",
X"44",
X"1B",
X"E5",
X"F1",
X"E9",
X"F0",
X"EB",
X"F1",
X"EC",
X"F1",
X"EC",
X"F0",
X"EB",
X"F4",
X"E6",
X"0A",
X"44",
X"3F",
X"3E",
X"42",
X"0C",
X"E4",
X"F2",
X"EA",
X"F1",
X"EB",
X"F1",
X"EC",
X"F1",
X"EC",
X"F2",
X"E9",
X"F4",
X"E7",
X"19",
X"48",
X"3F",
X"3E",
X"3F",
X"00",
X"E8",
X"F1",
X"EB",
X"F0",
X"EC",
X"EF",
X"EE",
X"F1",
X"EC",
X"F1",
X"EA",
X"F3",
X"EC",
X"28",
X"47",
X"3D",
X"41",
X"38",
X"F3",
X"ED",
X"F0",
X"ED",
X"EE",
X"ED",
X"F0",
X"F0",
X"EF",
X"EF",
X"EF",
X"EC",
X"EF",
X"F2",
X"34",
X"44",
X"3D",
X"43",
X"2C",
X"EE",
X"F0",
X"ED",
X"F1",
X"ED",
X"EF",
X"F0",
X"EF",
X"ED",
X"F2",
X"ED",
X"EE",
X"EC",
X"FC",
X"3C",
X"42",
X"40",
X"45",
X"20",
X"E8",
X"F4",
X"EC",
X"F2",
X"ED",
X"EF",
X"EE",
X"F2",
X"EA",
X"F5",
X"ED",
X"F1",
X"EB",
X"05",
X"42",
X"45",
X"3D",
X"42",
X"0D",
X"E8",
X"EF",
X"EE",
X"F3",
X"ED",
X"ED",
X"EE",
X"F3",
X"F2",
X"F0",
X"F7",
X"ED",
X"00",
X"41",
X"41",
X"41",
X"3F",
X"01",
X"E8",
X"F1",
X"EE",
X"EF",
X"EF",
X"EF",
X"EE",
X"F2",
X"ED",
X"F0",
X"F0",
X"EC",
X"24",
X"4E",
X"3D",
X"49",
X"24",
X"EF",
X"EC",
X"EF",
X"EF",
X"EE",
X"EC",
X"F0",
X"EC",
X"F3",
X"EC",
X"F0",
X"EA",
X"FA",
X"3D",
X"49",
X"41",
X"47",
X"08",
X"E6",
X"F0",
X"ED",
X"F2",
X"F1",
X"F0",
X"EE",
X"F0",
X"F0",
X"ED",
X"F0",
X"E8",
X"12",
X"4A",
X"3E",
X"46",
X"32",
X"F2",
X"EB",
X"EF",
X"ED",
X"F1",
X"F0",
X"F1",
X"F2",
X"F3",
X"EE",
X"EF",
X"EE",
X"F1",
X"31",
X"4A",
X"3B",
X"48",
X"16",
X"E7",
X"F0",
X"EE",
X"EF",
X"EF",
X"EE",
X"F2",
X"EF",
X"F1",
X"EE",
X"F3",
X"EB",
X"04",
X"3E",
X"38",
X"39",
X"37",
X"FC",
X"E9",
X"F0",
X"EE",
X"F1",
X"EF",
X"F2",
X"F1",
X"F0",
X"EE",
X"EF",
X"F3",
X"EC",
X"1E",
X"42",
X"31",
X"3F",
X"22",
X"EE",
X"F1",
X"F0",
X"EF",
X"F1",
X"F0",
X"F1",
X"F1",
X"F3",
X"ED",
X"F1",
X"ED",
X"FA",
X"36",
X"3B",
X"35",
X"3F",
X"06",
X"EA",
X"F3",
X"EF",
X"F2",
X"F0",
X"F2",
X"F1",
X"F0",
X"F0",
X"EE",
X"F4",
X"EC",
X"12",
X"43",
X"34",
X"3E",
X"2E",
X"F3",
X"EE",
X"F2",
X"EF",
X"F2",
X"F0",
X"F2",
X"EF",
X"F1",
X"EE",
X"F2",
X"F0",
X"F2",
X"2E",
X"3F",
X"32",
X"44",
X"13",
X"EB",
X"F3",
X"EF",
X"F1",
X"F2",
X"F2",
X"F1",
X"EF",
X"F0",
X"EE",
X"F3",
X"EC",
X"05",
X"40",
X"39",
X"3C",
X"39",
X"FB",
X"ED",
X"F3",
X"EE",
X"F2",
X"F1",
X"F0",
X"EE",
X"F4",
X"EF",
X"F0",
X"F4",
X"EE",
X"21",
X"42",
X"34",
X"42",
X"1E",
X"ED",
X"F3",
X"F1",
X"EF",
X"F2",
X"F0",
X"F0",
X"F0",
X"F2",
X"EF",
X"F7",
X"EE",
X"FF",
X"3C",
X"3B",
X"36",
X"3D",
X"03",
X"E7",
X"F4",
X"EF",
X"F0",
X"F2",
X"F2",
X"F2",
X"F3",
X"F3",
X"F1",
X"F4",
X"EE",
X"16",
X"44",
X"34",
X"3F",
X"29",
X"F1",
X"F0",
X"F0",
X"EF",
X"F3",
X"EC",
X"F1",
X"F2",
X"F2",
X"F2",
X"F5",
X"F1",
X"F6",
X"2F",
X"42",
X"34",
X"40",
X"0F",
X"E9",
X"F3",
X"ED",
X"F2",
X"F0",
X"F2",
X"F3",
X"F4",
X"F2",
X"F2",
X"F3",
X"F3",
X"2E",
X"3E",
X"32",
X"3A",
X"FE",
X"EC",
X"F3",
X"ED",
X"F3",
X"EE",
X"F1",
X"F1",
X"F4",
X"F3",
X"F4",
X"ED",
X"0F",
X"42",
X"34",
X"42",
X"1E",
X"EC",
X"F3",
X"EF",
X"F1",
X"F1",
X"F1",
X"F0",
X"F1",
X"F0",
X"F2",
X"F0",
X"F7",
X"35",
X"3C",
X"39",
X"38",
X"FB",
X"ED",
X"F2",
X"EF",
X"F4",
X"F3",
X"F4",
X"F2",
X"F5",
X"EF",
X"F3",
X"EF",
X"17",
X"41",
X"34",
X"3F",
X"16",
X"EB",
X"F4",
X"F0",
X"EF",
X"EF",
X"F2",
X"EF",
X"F4",
X"F4",
X"F5",
X"EF",
X"FD",
X"3D",
X"3C",
X"3B",
X"35",
X"F6",
X"EC",
X"F2",
X"F0",
X"EF",
X"EE",
X"F0",
X"F1",
X"F4",
X"F2",
X"F5",
X"ED",
X"1F",
X"43",
X"34",
X"40",
X"0F",
X"EB",
X"F5",
X"F2",
X"F2",
X"EC",
X"EF",
X"EE",
X"F1",
X"F0",
X"F5",
X"EF",
X"00",
X"41",
X"3A",
X"3B",
X"30",
X"F3",
X"F2",
X"F5",
X"F4",
X"F2",
X"EF",
X"F0",
X"EE",
X"EE",
X"EE",
X"F2",
X"EE",
X"26",
X"41",
X"32",
X"3F",
X"09",
X"EE",
X"F7",
X"F3",
X"F5",
X"EF",
X"F2",
X"EE",
X"EF",
X"EE",
X"F2",
X"EC",
X"03",
X"3B",
X"30",
X"38",
X"25",
X"EF",
X"F3",
X"F2",
X"F3",
X"F2",
X"F0",
X"F1",
X"EE",
X"EF",
X"EF",
X"F0",
X"F4",
X"2A",
X"3A",
X"2F",
X"36",
X"00",
X"EE",
X"F6",
X"F2",
X"F1",
X"ED",
X"F2",
X"F0",
X"F2",
X"F1",
X"F3",
X"ED",
X"0E",
X"3D",
X"2E",
X"38",
X"19",
X"EB",
X"F2",
X"F1",
X"F2",
X"F1",
X"F2",
X"F2",
X"F4",
X"F3",
X"F4",
X"F3",
X"F7",
X"2D",
X"34",
X"2C",
X"2F",
X"F9",
X"EF",
X"F5",
X"F0",
X"F6",
X"F1",
X"F3",
X"F4",
X"F3",
X"EF",
X"F7",
X"EF",
X"12",
X"3D",
X"28",
X"37",
X"13",
X"EB",
X"F7",
X"EE",
X"F2",
X"F0",
X"F0",
X"F4",
X"F7",
X"F3",
X"F3",
X"F0",
X"F7",
X"34",
X"36",
X"31",
X"31",
X"F6",
X"F0",
X"F4",
X"EE",
X"F3",
X"F0",
X"F3",
X"F6",
X"F4",
X"EF",
X"F6",
X"EA",
X"17",
X"40",
X"2D",
X"3E",
X"10",
X"EC",
X"F3",
X"ED",
X"F6",
X"F2",
X"F4",
X"F4",
X"F3",
X"EE",
X"F6",
X"EF",
X"FE",
X"36",
X"31",
X"36",
X"2A",
X"F6",
X"F2",
X"F1",
X"F2",
X"F3",
X"F3",
X"F3",
X"F4",
X"F1",
X"F2",
X"F4",
X"F9",
X"32",
X"33",
X"35",
X"26",
X"F3",
X"F3",
X"F0",
X"F1",
X"F2",
X"F3",
X"F2",
X"F4",
X"EE",
X"F3",
X"F4",
X"1A",
X"3C",
X"2F",
X"34",
X"00",
X"EF",
X"F5",
X"F0",
X"F5",
X"F3",
X"F3",
X"F3",
X"F0",
X"F2",
X"F1",
X"02",
X"39",
X"31",
X"37",
X"18",
X"EC",
X"F4",
X"F0",
X"F3",
X"F4",
X"F4",
X"F3",
X"F4",
X"F1",
X"F3",
X"F3",
X"2A",
X"37",
X"32",
X"2F",
X"F4",
X"F1",
X"F1",
X"F1",
X"F2",
X"F3",
X"F2",
X"F3",
X"F1",
X"F5",
X"F0",
X"12",
X"3C",
X"2E",
X"39",
X"07",
X"EC",
X"F4",
X"F0",
X"F2",
X"F4",
X"F3",
X"F3",
X"F3",
X"F2",
X"F1",
X"FD",
X"36",
X"32",
X"38",
X"20",
X"EE",
X"F3",
X"F0",
X"F2",
X"F2",
X"F4",
X"F1",
X"F4",
X"F0",
X"F4",
X"F0",
X"20",
X"38",
X"30",
X"35",
X"FB",
X"EF",
X"F3",
X"F2",
X"F3",
X"F4",
X"F1",
X"F3",
X"F1",
X"F4",
X"EF",
X"07",
X"3A",
X"2D",
X"3A",
X"0F",
X"EB",
X"F4",
X"F1",
X"F4",
X"F3",
X"F3",
X"F1",
X"F2",
X"F2",
X"F3",
X"F4",
X"2F",
X"33",
X"35",
X"29",
X"F1",
X"F3",
X"F3",
X"F4",
X"F2",
X"F2",
X"F1",
X"F4",
X"F1",
X"F6",
X"ED",
X"18",
X"3C",
X"2E",
X"38",
X"00",
X"EF",
X"F4",
X"F2",
X"F2",
X"F2",
X"F2",
X"F3",
X"F2",
X"F3",
X"EF",
X"00",
X"3A",
X"30",
X"39",
X"18",
X"ED",
X"F6",
X"F0",
X"F3",
X"F1",
X"F3",
X"F2",
X"F3",
X"F0",
X"F3",
X"F1",
X"23",
X"30",
X"2C",
X"28",
X"F4",
X"F1",
X"F0",
X"F3",
X"F3",
X"F3",
X"F2",
X"F1",
X"F0",
X"F4",
X"EF",
X"0C",
X"35",
X"28",
X"33",
X"06",
X"ED",
X"F2",
X"F1",
X"F3",
X"F2",
X"F3",
X"F1",
X"F3",
X"F3",
X"F3",
X"F9",
X"2D",
X"2A",
X"30",
X"1C",
X"F0",
X"F4",
X"F1",
X"F3",
X"F0",
X"F4",
X"F1",
X"F3",
X"F2",
X"F5",
X"F0",
X"1C",
X"31",
X"2A",
X"2F",
X"FB",
X"F1",
X"F1",
X"F2",
X"F3",
X"F3",
X"F3",
X"F3",
X"F2",
X"F4",
X"F0",
X"05",
X"34",
X"26",
X"34",
X"0D",
X"EE",
X"F4",
X"EF",
X"F3",
X"F2",
X"F6",
X"F3",
X"F4",
X"F2",
X"F3",
X"F6",
X"28",
X"2D",
X"2E",
X"24",
X"F1",
X"F3",
X"F0",
X"F4",
X"F3",
X"F5",
X"F2",
X"F5",
X"F1",
X"F4",
X"EF",
X"15",
X"30",
X"2A",
X"2B",
X"F5",
X"F5",
X"F2",
X"F2",
X"F3",
X"F2",
X"F4",
X"F4",
X"F4",
X"F2",
X"00",
X"31",
X"28",
X"31",
X"04",
X"EE",
X"F4",
X"F3",
X"F2",
X"F4",
X"F2",
X"F4",
X"F3",
X"F6",
X"F3",
X"24",
X"2E",
X"2E",
X"1D",
X"EE",
X"F5",
X"F1",
X"F4",
X"F1",
X"F2",
X"F3",
X"F3",
X"F6",
X"F0",
X"0D",
X"35",
X"28",
X"2F",
X"F9",
X"F2",
X"F1",
X"F3",
X"F0",
X"F5",
X"F2",
X"F6",
X"F3",
X"F4",
X"FA",
X"2F",
X"28",
X"33",
X"0E",
X"EF",
X"F4",
X"F1",
X"F2",
X"F2",
X"F3",
X"F3",
X"F3",
X"F5",
X"F0",
X"1C",
X"31",
X"2C",
X"26",
X"F1",
X"F4",
X"F1",
X"F3",
X"F2",
X"F3",
X"F2",
X"F2",
X"F4",
X"F1",
X"04",
X"35",
X"28",
X"33",
X"00",
X"F0",
X"F3",
X"F3",
X"F3",
X"F4",
X"F2",
X"F5",
X"F3",
X"F4",
X"F5",
X"2A",
X"2C",
X"32",
X"16",
X"ED",
X"F5",
X"F2",
X"F2",
X"F3",
X"F4",
X"F5",
X"F3",
X"F6",
X"EF",
X"14",
X"34",
X"2A",
X"2A",
X"F6",
X"F3",
X"F2",
X"F4",
X"F1",
X"F4",
X"F3",
X"F5",
X"F5",
X"F2",
X"FF",
X"32",
X"28",
X"34",
X"06",
X"EF",
X"F4",
X"F2",
X"F3",
X"F3",
X"F3",
X"F4",
X"F2",
X"F5",
X"F1",
X"24",
X"2E",
X"2F",
X"1F",
X"EF",
X"F5",
X"F1",
X"F3",
X"F2",
X"F4",
X"F4",
X"F2",
X"F5",
X"EE",
X"0C",
X"34",
X"29",
X"30",
X"FA",
X"F3",
X"F3",
X"F3",
X"F2",
X"F3",
X"F2",
X"F4",
X"F3",
X"F3",
X"F9",
X"2F",
X"2A",
X"34",
X"0F",
X"EF",
X"F4",
X"F2",
X"F2",
X"F2",
X"F3",
X"F3",
X"F4",
X"F7",
X"EF",
X"1C",
X"31",
X"2D",
X"27",
X"F1",
X"F3",
X"F2",
X"F4",
X"F1",
X"F4",
X"F2",
X"F4",
X"F5",
X"F1",
X"00",
X"2C",
X"20",
X"2C",
X"00",
X"F1",
X"F3",
X"F3",
X"F2",
X"F4",
X"F1",
X"F5",
X"F4",
X"F5",
X"F5",
X"22",
X"25",
X"2A",
X"14",
X"EF",
X"F5",
X"F2",
X"F3",
X"F4",
X"F1",
X"F4",
X"F3",
X"F5",
X"F1",
X"0F",
X"2A",
X"26",
X"26",
X"F7",
X"F5",
X"F2",
X"F2",
X"F3",
X"F2",
X"F5",
X"F3",
X"F5",
X"F2",
X"FE",
X"2A",
X"22",
X"2C",
X"06",
X"F1",
X"F4",
X"F2",
X"F0",
X"F3",
X"F3",
X"F5",
X"F4",
X"F5",
X"F3",
X"1D",
X"27",
X"28",
X"1A",
X"F1",
X"F8",
X"F2",
X"F2",
X"F2",
X"F2",
X"F4",
X"F6",
X"F4",
X"F6",
X"21",
X"25",
X"27",
X"09",
X"ED",
X"F9",
X"F0",
X"F7",
X"F2",
X"F8",
X"F1",
X"F8",
X"EE",
X"0C",
X"2A",
X"25",
X"1E",
X"F3",
X"F4",
X"F4",
X"F4",
X"F4",
X"F4",
X"F5",
X"F6",
X"F3",
X"FA",
X"24",
X"24",
X"29",
X"03",
X"EF",
X"F7",
X"F1",
X"F6",
X"F4",
X"F7",
X"F2",
X"F8",
X"F0",
X"13",
X"29",
X"25",
X"1C",
X"F1",
X"F5",
X"F2",
X"F6",
X"F3",
X"F6",
X"F3",
X"F6",
X"F3",
X"FE",
X"26",
X"26",
X"27",
X"00",
X"EF",
X"F6",
X"F2",
X"F7",
X"F3",
X"F7",
X"F2",
X"F8",
X"F0",
X"18",
X"27",
X"27",
X"16",
X"EF",
X"F7",
X"F2",
X"F7",
X"F3",
X"F8",
X"F3",
X"F7",
X"F1",
X"01",
X"29",
X"25",
X"25",
X"FB",
X"F2",
X"F6",
X"F4",
X"F6",
X"F4",
X"F6",
X"F3",
X"F7",
X"F2",
X"1D",
X"27",
X"28",
X"10",
X"EF",
X"F8",
X"F2",
X"F7",
X"F2",
X"F8",
X"F2",
X"F8",
X"F0",
X"07",
X"29",
X"25",
X"24",
X"F7",
X"F4",
X"F4",
X"F4",
X"F5",
X"F4",
X"F5",
X"F4",
X"F6",
X"F5",
X"22",
X"26",
X"29",
X"0B",
X"EF",
X"F8",
X"F1",
X"F8",
X"F2",
X"F7",
X"F2",
X"F9",
X"F0",
X"0D",
X"2A",
X"26",
X"20",
X"F3",
X"F5",
X"F3",
X"F5",
X"F4",
X"F6",
X"F4",
X"F5",
X"F4",
X"F9",
X"25",
X"25",
X"29",
X"04",
X"F0",
X"F7",
X"F2",
X"F8",
X"F3",
X"F7",
X"F1",
X"F9",
X"EF",
X"13",
X"29",
X"27",
X"1B",
X"F0",
X"F6",
X"F2",
X"F6",
X"F4",
X"F6",
X"F4",
X"F6",
X"F3",
X"FD",
X"27",
X"25",
X"28",
X"00",
X"F0",
X"F7",
X"F3",
X"F7",
X"F3",
X"F7",
X"F2",
X"F8",
X"F0",
X"18",
X"28",
X"28",
X"16",
X"EF",
X"F7",
X"F2",
X"F7",
X"F3",
X"F7",
X"F3",
X"F7",
X"F0",
X"00",
X"29",
X"25",
X"27",
X"FC",
X"F2",
X"F6",
X"F3",
X"F7",
X"F4",
X"F6",
X"F3",
X"F7",
X"F1",
X"1D",
X"27",
X"29",
X"11",
X"EE",
X"F7",
X"F1",
X"F7",
X"F4",
X"F7",
X"F2",
X"F8",
X"F1",
X"03",
X"21",
X"1E",
X"1D",
X"F8",
X"F4",
X"F6",
X"F5",
X"F5",
X"F4",
X"F5",
X"F5",
X"F6",
X"F6",
X"1A",
X"1E",
X"21",
X"08",
X"F1",
X"F9",
X"F2",
X"F6",
X"F2",
X"F7",
X"F3",
X"F8",
X"F2",
X"08",
X"22",
X"1E",
X"1A",
X"F5",
X"F7",
X"F4",
X"F5",
X"F2",
X"F7",
X"F2",
X"F9",
X"F1",
X"0C",
X"21",
X"20",
X"0F",
X"F2",
X"F8",
X"F3",
X"F8",
X"F4",
X"F7",
X"F3",
X"F5",
X"F7",
X"1D",
X"1F",
X"20",
X"FE",
X"F4",
X"F6",
X"F5",
X"F4",
X"F7",
X"F4",
X"F9",
X"F2",
X"05",
X"23",
X"1F",
X"16",
X"F3",
X"F8",
X"F4",
X"F7",
X"F3",
X"F7",
X"F3",
X"F8",
X"F3",
X"17",
X"21",
X"21",
X"04",
X"F3",
X"F7",
X"F5",
X"F4",
X"F4",
X"F6",
X"F7",
X"F5",
X"FF",
X"22",
X"1F",
X"1C",
X"F5",
X"F8",
X"F4",
X"F7",
X"F2",
X"F7",
X"F4",
X"FA",
X"F2",
X"10",
X"22",
X"22",
X"0D",
X"F0",
X"F8",
X"F3",
X"F7",
X"F4",
X"F7",
X"F6",
X"F7",
X"FA",
X"1E",
X"1F",
X"20",
X"FC",
X"F5",
X"F5",
X"F7",
X"F5",
X"F8",
X"F4",
X"FA",
X"F1",
X"09",
X"21",
X"21",
X"14",
X"F1",
X"F9",
X"F3",
X"F9",
X"F4",
X"F8",
X"F4",
X"F8",
X"F4",
X"1A",
X"1F",
X"22",
X"01",
X"F2",
X"F8",
X"F5",
X"F7",
X"F6",
X"F6",
X"F8",
X"F4",
X"00",
X"22",
X"1F",
X"1A",
X"F4",
X"F8",
X"F4",
X"F8",
X"F4",
X"F8",
X"F4",
X"FA",
X"F2",
X"14",
X"20",
X"22",
X"09",
X"F2",
X"F8",
X"F5",
X"F7",
X"F5",
X"F6",
X"F6",
X"F6",
X"FB",
X"20",
X"1E",
X"20",
X"F9",
X"F6",
X"F5",
X"F8",
X"F5",
X"F8",
X"F4",
X"FA",
X"F2",
X"0C",
X"21",
X"21",
X"11",
X"F1",
X"F9",
X"F4",
X"F8",
X"F4",
X"F7",
X"F5",
X"F8",
X"F7",
X"1C",
X"1F",
X"21",
X"00",
X"F4",
X"F7",
X"F7",
X"F6",
X"F7",
X"F5",
X"F8",
X"F3",
X"04",
X"22",
X"1F",
X"19",
X"F3",
X"F9",
X"F4",
X"F8",
X"F4",
X"F8",
X"F5",
X"FA",
X"F3",
X"17",
X"1F",
X"23",
X"06",
X"F3",
X"F8",
X"F4",
X"F7",
X"F5",
X"F7",
X"F7",
X"F6",
X"FF",
X"22",
X"1F",
X"1F",
X"F7",
X"F7",
X"F4",
X"F7",
X"F5",
X"F8",
X"F4",
X"FB",
X"F2",
X"0F",
X"22",
X"22",
X"0F",
X"F1",
X"FA",
X"F3",
X"F9",
X"F4",
X"F8",
X"F5",
X"F9",
X"F8",
X"1F",
X"1E",
X"22",
X"FD",
X"F6",
X"F5",
X"F7",
X"F5",
X"F8",
X"F5",
X"FA",
X"F2",
X"07",
X"23",
X"21",
X"17",
X"F1",
X"F9",
X"F4",
X"F7",
X"F4",
X"F9",
X"F5",
X"F9",
X"F3",
X"1A",
X"20",
X"22",
X"02",
X"F2",
X"F8",
X"F5",
X"F8",
X"F7",
X"F6",
X"F7",
X"F3",
X"0A",
X"1A",
X"18",
X"01",
X"F2",
X"F9",
X"F5",
X"F9",
X"F6",
X"F8",
X"F6",
X"F7",
X"10",
X"1A",
X"15",
X"FE",
X"F3",
X"FA",
X"F4",
X"FA",
X"F5",
X"F9",
X"F4",
X"FB",
X"14",
X"1A",
X"12",
X"FA",
X"F5",
X"F9",
X"F5",
X"F9",
X"F5",
X"FA",
X"F3",
X"00",
X"17",
X"1B",
X"0E",
X"F6",
X"F8",
X"F8",
X"F6",
X"F9",
X"F6",
X"FA",
X"F3",
X"05",
X"1A",
X"1A",
X"08",
X"F4",
X"F9",
X"F7",
X"F7",
X"F7",
X"F7",
X"F9",
X"F4",
X"0B",
X"1A",
X"19",
X"02",
X"F3",
X"FA",
X"F6",
X"F9",
X"F7",
X"F8",
X"F8",
X"F8",
X"11",
X"1B",
X"17",
X"FE",
X"F4",
X"FA",
X"F5",
X"F9",
X"F5",
X"FA",
X"F6",
X"FC",
X"15",
X"1B",
X"13",
X"FA",
X"F6",
X"F9",
X"F6",
X"F9",
X"F6",
X"FA",
X"F4",
X"00",
X"18",
X"1B",
X"0F",
X"F6",
X"F7",
X"F8",
X"F7",
X"F9",
X"F6",
X"FA",
X"F4",
X"05",
X"1A",
X"1B",
X"0A",
X"F4",
X"F9",
X"F6",
X"F8",
X"F8",
X"F7",
X"F9",
X"F5",
X"0C",
X"1B",
X"19",
X"04",
X"F4",
X"FA",
X"F6",
X"F9",
X"F6",
X"F9",
X"F8",
X"F8",
X"11",
X"1C",
X"17",
X"FF",
X"F4",
X"FA",
X"F6",
X"FA",
X"F6",
X"FA",
X"F6",
X"FD",
X"16",
X"1C",
X"14",
X"FA",
X"F6",
X"F9",
X"F6",
X"FA",
X"F6",
X"FB",
X"F5",
X"01",
X"19",
X"1B",
X"0F",
X"F7",
X"F8",
X"F8",
X"F7",
X"F9",
X"F6",
X"FA",
X"F5",
X"06",
X"1A",
X"1B",
X"0A",
X"F5",
X"FA",
X"F7",
X"F9",
X"F8",
X"F8",
X"F9",
X"F5",
X"0C",
X"1C",
X"19",
X"04",
X"F4",
X"FB",
X"F7",
X"FA",
X"F7",
X"F9",
X"F8",
X"F8",
X"11",
X"1C",
X"17",
X"00",
X"F5",
X"FB",
X"F6",
X"FA",
X"F6",
X"FA",
X"F6",
X"FD",
X"15",
X"1C",
X"14",
X"FB",
X"F6",
X"FA",
X"F7",
X"FA",
X"F6",
X"FB",
X"F5",
X"00",
X"19",
X"1C",
X"0F",
X"F7",
X"F8",
X"F9",
X"F8",
X"FA",
X"F6",
X"FB",
X"F4",
X"07",
X"1B",
X"1B",
X"0A",
X"F5",
X"FA",
X"F8",
X"F8",
X"F9",
X"F8",
X"FA",
X"F5",
X"0D",
X"1C",
X"1A",
X"04",
X"F4",
X"FA",
X"F7",
X"FA",
X"F8",
X"F8",
X"F8",
X"F8",
X"12",
X"1D",
X"18",
X"00",
X"F4",
X"FA",
X"F7",
X"FB",
X"F7",
X"FA",
X"F7",
X"FD",
X"16",
X"1E",
X"0F",
X"F7",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F8",
X"FC",
X"16",
X"1C",
X"11",
X"F6",
X"F9",
X"F7",
X"F9",
X"F7",
X"FA",
X"F8",
X"FC",
X"15",
X"1D",
X"10",
X"F7",
X"F9",
X"F8",
X"F9",
X"F8",
X"F8",
X"F8",
X"FA",
X"0E",
X"13",
X"0B",
X"F7",
X"F9",
X"F8",
X"FA",
X"F8",
X"F9",
X"F8",
X"FB",
X"0D",
X"13",
X"0B",
X"F8",
X"F9",
X"F8",
X"F9",
X"F9",
X"F9",
X"F8",
X"FA",
X"0E",
X"13",
X"0C",
X"F8",
X"F9",
X"F8",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"0D",
X"13",
X"0C",
X"F8",
X"F9",
X"F9",
X"FA",
X"F9",
X"F9",
X"F9",
X"FA",
X"0D",
X"13",
X"0D",
X"F9",
X"F9",
X"F9",
X"FA",
X"F9",
X"F9",
X"F9",
X"FA",
X"0E",
X"13",
X"0D",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"0E",
X"14",
X"0D",
X"F9",
X"F9",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"0D",
X"14",
X"0E",
X"FA",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FA",
X"0D",
X"14",
X"0E",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"F9",
X"FA",
X"F9",
X"0E",
X"14",
X"0E",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"F9",
X"FA",
X"FA",
X"0D",
X"15",
X"0F",
X"FB",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"F9",
X"0D",
X"15",
X"0F",
X"FB",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FB",
X"F9",
X"0D",
X"15",
X"0F",
X"FC",
X"F9",
X"FA",
X"F9",
X"FB",
X"F9",
X"FB",
X"F9",
X"0D",
X"15",
X"10",
X"FC",
X"F9",
X"FA",
X"F9",
X"FB",
X"F9",
X"FB",
X"F9",
X"0D",
X"14",
X"10",
X"FC",
X"F9",
X"FB",
X"F9",
X"FB",
X"F9",
X"FB",
X"F9",
X"0C",
X"14",
X"10",
X"FD",
X"FA",
X"FB",
X"FA",
X"FB",
X"F9",
X"FB",
X"F9",
X"0C",
X"14",
X"10",
X"FD",
X"FA",
X"FB",
X"F9",
X"FB",
X"F9",
X"FB",
X"F8",
X"0C",
X"15",
X"10",
X"FD",
X"F9",
X"FB",
X"F9",
X"FB",
X"FA",
X"FC",
X"F9",
X"0B",
X"15",
X"10",
X"FD",
X"F9",
X"FB",
X"F9",
X"FB",
X"FA",
X"FC",
X"F9",
X"0C",
X"14",
X"11",
X"FE",
X"F9",
X"FB",
X"FA",
X"FB",
X"FA",
X"FC",
X"F9",
X"0B",
X"15",
X"11",
X"FE",
X"F9",
X"FB",
X"F9",
X"FB",
X"F9",
X"FC",
X"F8",
X"0B",
X"15",
X"11",
X"FE",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"F9",
X"00",
X"13",
X"14",
X"03",
X"F8",
X"FC",
X"F9",
X"FB",
X"FA",
X"FB",
X"FB",
X"0F",
X"15",
X"0A",
X"F8",
X"FC",
X"F9",
X"FC",
X"F9",
X"FD",
X"F8",
X"09",
X"15",
X"10",
X"FB",
X"FA",
X"FA",
X"FB",
X"FA",
X"FC",
X"F8",
X"02",
X"14",
X"13",
X"00",
X"F8",
X"FC",
X"F9",
X"FB",
X"FA",
X"FB",
X"FD",
X"11",
X"15",
X"08",
X"F7",
X"FC",
X"F9",
X"FC",
X"F9",
X"FC",
X"F9",
X"0C",
X"15",
X"0F",
X"FA",
X"FB",
X"F9",
X"FC",
X"FA",
X"FC",
X"F9",
X"01",
X"0C",
X"0B",
X"FE",
X"FA",
X"FB",
X"FA",
X"FA",
X"FB",
X"FA",
X"FE",
X"0B",
X"0C",
X"02",
X"F8",
X"FC",
X"FA",
X"FC",
X"FA",
X"FC",
X"FA",
X"08",
X"0D",
X"07",
X"F9",
X"FC",
X"FA",
X"FC",
X"FA",
X"FC",
X"F9",
X"03",
X"0D",
X"0A",
X"FD",
X"FA",
X"FB",
X"FB",
X"FB",
X"FC",
X"FA",
X"00",
X"0B",
X"0C",
X"00",
X"F9",
X"FC",
X"FA",
X"FC",
X"FB",
X"FC",
X"FC",
X"09",
X"0C",
X"05",
X"F9",
X"FD",
X"FA",
X"FD",
X"FA",
X"FD",
X"FA",
X"05",
X"0D",
X"09",
X"FC",
X"FC",
X"FB",
X"FC",
X"FB",
X"FD",
X"FA",
X"00",
X"0C",
X"0C",
X"00",
X"FA",
X"FC",
X"FB",
X"FC",
X"FB",
X"FB",
X"FD",
X"0A",
X"0D",
X"04",
X"F9",
X"FD",
X"FB",
X"FD",
X"FB",
X"FD",
X"FA",
X"07",
X"0D",
X"09",
X"FB",
X"FC",
X"FB",
X"FD",
X"FB",
X"FD",
X"FA",
X"02",
X"0D",
X"0C",
X"FF",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FB",
X"FF",
X"0C",
X"0D",
X"02",
X"FA",
X"FD",
X"FB",
X"FD",
X"FB",
X"FD",
X"FB",
X"09",
X"0D",
X"07",
X"FB",
X"FD",
X"FB",
X"FD",
X"FB",
X"FD",
X"FA",
X"04",
X"0D",
X"0B",
X"FE",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FB",
X"00",
X"0C",
X"0D",
X"01",
X"FA",
X"FD",
X"FB",
X"FD",
X"FC",
X"FD",
X"FD",
X"0A",
X"0D",
X"06",
X"FA",
X"FE",
X"FB",
X"FD",
X"FB",
X"FE",
X"FA",
X"06",
X"0D",
X"0A",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FE",
X"FA",
X"01",
X"0D",
X"0D",
X"00",
X"FB",
X"FD",
X"FC",
X"FD",
X"FD",
X"FC",
X"FF",
X"0B",
X"0D",
X"04",
X"FA",
X"FD",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"07",
X"0F",
X"06",
X"FB",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FF",
X"0B",
X"0E",
X"01",
X"FB",
X"FD",
X"FC",
X"FD",
X"FD",
X"FC",
X"02",
X"0F",
X"0A",
X"FE",
X"FB",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"07",
X"0F",
X"05",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"00",
X"0C",
X"0E",
X"00",
X"FB",
X"FD",
X"FD",
X"FD",
X"FD",
X"FB",
X"02",
X"0F",
X"0A",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"08",
X"10",
X"04",
X"FB",
X"FD",
X"FD",
X"FC",
X"FD",
X"FB",
X"00",
X"0C",
X"0E",
X"00",
X"FB",
X"FD",
X"FC",
X"FD",
X"FD",
X"FC",
X"03",
X"0F",
X"09",
X"FE",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"08",
X"0F",
X"04",
X"FC",
X"FD",
X"FD",
X"FC",
X"FD",
X"FB",
X"00",
X"0D",
X"0D",
X"00",
X"FB",
X"FD",
X"FC",
X"FD",
X"FD",
X"FC",
X"00",
X"05",
X"02",
X"FD",
X"FD",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"02",
X"05",
X"00",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FC",
X"FF",
X"04",
X"04",
X"FF",
X"FD",
X"FE",
X"FD",
X"FD",
X"FD",
X"FD",
X"00",
X"05",
X"02",
X"FD",
X"FD",
X"FE",
X"FD",
X"FD",
X"FD",
X"FE",
X"03",
X"06",
X"00",
X"FD",
X"FE",
X"FD",
X"FD",
X"FE",
X"FD",
X"00",
X"05",
X"04",
X"FF",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FD",
X"01",
X"06",
X"02",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"03",
X"06",
X"00",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FD",
X"00",
X"05",
X"04",
X"00",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"01",
X"06",
X"02",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FD",
X"FF",
X"04",
X"06",
X"00",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"00",
X"06",
X"04",
X"FF",
X"FE",
X"FF",
X"FE",
X"FE",
X"FE",
X"FE",
X"02",
X"06",
X"02",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"04",
X"06",
X"00",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"00",
X"06",
X"04",
X"00",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF" );
--//--------------------------------------
  begin

    if (RESET_N='0') then
      Q <= sqr_table(0);
    elsif(rising_edge(CLK)) then
      if (ENA='1') then
          Q <= sqr_table(to_integer(unsigned(ADDR)));
      end if;
    end if;
  end process;
end arch;