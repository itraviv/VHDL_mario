--------------------------------------
-- SinTable.vhd
-- Written by Saar Eliad and Itamar Raviv.
-- All rights reserved, Copyright 2017
--------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ThemeSoundTable is
port(
  CLK     : in std_logic;
  RESET_N : in std_logic;
  ENA     : in std_logic;
  ADDR    : in std_logic_vector(11 downto 0);
  Q       : out std_logic_vector(7 downto 0)
);
end ThemeSoundTable;

architecture arch of ThemeSoundTable is

type table_type is array(0 to 4095) of std_logic_vector(7 downto 0);
signal sqr_table : table_type;

begin

  SQRTableTC_proc: process(RESET_N, CLK)
    constant sqr_table : table_type := (
	X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FE",
X"00",
X"FF",
X"01",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"02",
X"FD",
X"01",
X"FF",
X"00",
X"00",
X"02",
X"FA",
X"02",
X"FC",
X"03",
X"FB",
X"04",
X"FE",
X"07",
X"F8",
X"07",
X"F4",
X"10",
X"F9",
X"2C",
X"5A",
X"56",
X"4F",
X"4E",
X"4F",
X"37",
X"39",
X"2F",
X"38",
X"23",
X"2C",
X"1D",
X"3A",
X"0B",
X"0D",
X"09",
X"07",
X"06",
X"00",
X"01",
X"00",
X"00",
X"EA",
X"F7",
X"F2",
X"F7",
X"F2",
X"F7",
X"09",
X"14",
X"E9",
X"FC",
X"FC",
X"FE",
X"00",
X"09",
X"11",
X"0A",
X"1B",
X"0F",
X"2B",
X"11",
X"25",
X"19",
X"33",
X"22",
X"3F",
X"2E",
X"2C",
X"34",
X"27",
X"36",
X"39",
X"3B",
X"35",
X"34",
X"36",
X"24",
X"1A",
X"17",
X"0E",
X"14",
X"18",
X"1B",
X"F0",
X"F0",
X"F1",
X"E9",
X"00",
X"DB",
X"E2",
X"D8",
X"E8",
X"D7",
X"E1",
X"D6",
X"EA",
X"D5",
X"D0",
X"D2",
X"DF",
X"E0",
X"D8",
X"E7",
X"F9",
X"FB",
X"EF",
X"E7",
X"F5",
X"FF",
X"FB",
X"FF",
X"07",
X"11",
X"16",
X"15",
X"13",
X"35",
X"12",
X"10",
X"24",
X"1A",
X"2E",
X"1E",
X"2E",
X"26",
X"27",
X"2A",
X"35",
X"29",
X"24",
X"24",
X"1D",
X"1E",
X"10",
X"14",
X"0B",
X"04",
X"01",
X"0C",
X"F3",
X"F2",
X"EF",
X"EB",
X"E1",
X"F8",
X"E2",
X"E9",
X"D4",
X"09",
X"0F",
X"1C",
X"25",
X"17",
X"0E",
X"15",
X"1C",
X"14",
X"E7",
X"D4",
X"E2",
X"F4",
X"BD",
X"F1",
X"05",
X"14",
X"0F",
X"14",
X"1C",
X"24",
X"22",
X"1E",
X"31",
X"22",
X"34",
X"27",
X"65",
X"60",
X"6A",
X"62",
X"42",
X"34",
X"0C",
X"03",
X"00",
X"00",
X"FD",
X"ED",
X"20",
X"21",
X"08",
X"34",
X"35",
X"37",
X"10",
X"0E",
X"EC",
X"E2",
X"E4",
X"DC",
X"03",
X"0C",
X"EF",
X"CD",
X"E3",
X"DA",
X"B3",
X"99",
X"B1",
X"A9",
X"C1",
X"A5",
X"E2",
X"2D",
X"18",
X"23",
X"26",
X"2C",
X"1C",
X"09",
X"09",
X"FE",
X"05",
X"FE",
X"00",
X"1F",
X"18",
X"14",
X"1D",
X"36",
X"08",
X"E4",
X"01",
X"F1",
X"18",
X"26",
X"42",
X"5A",
X"60",
X"4B",
X"4D",
X"4A",
X"2B",
X"02",
X"0E",
X"F4",
X"CC",
X"C7",
X"D1",
X"FB",
X"F1",
X"F9",
X"EC",
X"EB",
X"E6",
X"B5",
X"DB",
X"EF",
X"DA",
X"E2",
X"E1",
X"05",
X"08",
X"10",
X"F8",
X"FA",
X"0D",
X"AB",
X"AB",
X"C5",
X"BA",
X"C8",
X"C1",
X"00",
X"16",
X"08",
X"0E",
X"1C",
X"3C",
X"25",
X"15",
X"1C",
X"0C",
X"2B",
X"13",
X"3C",
X"57",
X"54",
X"2C",
X"25",
X"20",
X"FC",
X"EE",
X"EE",
X"E2",
X"E8",
X"E9",
X"FF",
X"0F",
X"0B",
X"39",
X"25",
X"21",
X"0B",
X"E4",
X"F9",
X"F7",
X"F4",
X"CC",
X"E7",
X"E9",
X"CD",
X"E0",
X"C9",
X"D2",
X"C5",
X"B7",
X"9B",
X"A5",
X"AF",
X"B8",
X"E9",
X"07",
X"16",
X"1C",
X"18",
X"1D",
X"15",
X"0B",
X"0C",
X"FA",
X"0C",
X"F3",
X"F0",
X"12",
X"0B",
X"1F",
X"17",
X"2B",
X"20",
X"0A",
X"09",
X"F9",
X"23",
X"3B",
X"20",
X"52",
X"45",
X"54",
X"3F",
X"43",
X"31",
X"1B",
X"F8",
X"D8",
X"E1",
X"D8",
X"CB",
X"E8",
X"F0",
X"F4",
X"F6",
X"FF",
X"E0",
X"D4",
X"DB",
X"D8",
X"E0",
X"DF",
X"DD",
X"DC",
X"00",
X"F8",
X"FF",
X"00",
X"00",
X"D9",
X"B6",
X"AB",
X"C6",
X"CA",
X"C9",
X"D9",
X"04",
X"04",
X"14",
X"26",
X"34",
X"43",
X"0D",
X"0D",
X"1C",
X"16",
X"2E",
X"20",
X"44",
X"54",
X"1E",
X"1C",
X"28",
X"25",
X"03",
X"F4",
X"FF",
X"00",
X"EF",
X"F1",
X"11",
X"28",
X"37",
X"33",
X"2E",
X"11",
X"FE",
X"E8",
X"EB",
X"ED",
X"DD",
X"D7",
X"D6",
X"DD",
X"DA",
X"DC",
X"D7",
X"CE",
X"B9",
X"A2",
X"B9",
X"B4",
X"C7",
X"E4",
X"FA",
X"1B",
X"13",
X"05",
X"1B",
X"20",
X"04",
X"F8",
X"05",
X"F5",
X"EB",
X"FC",
X"FD",
X"14",
X"1B",
X"0A",
X"14",
X"18",
X"1D",
X"FD",
X"1A",
X"32",
X"3D",
X"25",
X"35",
X"4D",
X"3B",
X"3A",
X"27",
X"3A",
X"20",
X"EC",
X"DC",
X"DC",
X"E6",
X"DD",
X"D4",
X"00",
X"E0",
X"EC",
X"E9",
X"EB",
X"00",
X"DF",
X"E7",
X"E5",
X"D1",
X"D3",
X"DF",
X"F1",
X"00",
X"F9",
X"EB",
X"D8",
X"DF",
X"C7",
X"D3",
X"CA",
X"D0",
X"DF",
X"DB",
X"07",
X"19",
X"14",
X"29",
X"26",
X"2F",
X"22",
X"1D",
X"0B",
X"13",
X"1E",
X"20",
X"42",
X"2E",
X"22",
X"2D",
X"2D",
X"21",
X"16",
X"0D",
X"FC",
X"E5",
X"FC",
X"DB",
X"1F",
X"30",
X"16",
X"1B",
X"17",
X"16",
X"08",
X"EE",
X"E5",
X"EF",
X"E6",
X"C7",
X"D2",
X"DB",
X"D9",
X"E9",
X"DA",
X"E7",
X"CC",
X"B2",
X"B0",
X"B3",
X"E1",
X"ED",
X"FB",
X"0F",
X"14",
X"1C",
X"10",
X"27",
X"27",
X"EE",
X"FA",
X"DA",
X"E7",
X"EE",
X"FB",
X"0F",
X"0D",
X"16",
X"1B",
X"2C",
X"1F",
X"0A",
X"33",
X"28",
X"25",
X"3C",
X"31",
X"1E",
X"37",
X"1D",
X"2B",
X"19",
X"10",
X"EB",
X"D8",
X"DB",
X"D2",
X"D8",
X"D2",
X"EF",
X"E9",
X"F8",
X"ED",
X"00",
X"FC",
X"E5",
X"DB",
X"DF",
X"E3",
X"E8",
X"DA",
X"E0",
X"F3",
X"E0",
X"DC",
X"D7",
X"E6",
X"D8",
X"CD",
X"E0",
X"F0",
X"D1",
X"E0",
X"F1",
X"FD",
X"1D",
X"22",
X"2F",
X"27",
X"2B",
X"11",
X"2B",
X"07",
X"26",
X"1E",
X"27",
X"28",
X"26",
X"38",
X"35",
X"23",
X"1D",
X"FB",
X"03",
X"FA",
X"F7",
X"FF",
X"17",
X"3A",
X"1D",
X"16",
X"18",
X"12",
X"0C",
X"00",
X"D7",
X"E6",
X"DD",
X"C4",
X"C5",
X"D4",
X"DF",
X"D9",
X"E0",
X"D6",
X"DE",
X"C6",
X"AF",
X"C8",
X"E5",
X"E5",
X"E7",
X"05",
X"1C",
X"04",
X"13",
X"16",
X"18",
X"10",
X"EE",
X"EB",
X"E6",
X"F4",
X"FD",
X"09",
X"1B",
X"1C",
X"29",
X"31",
X"37",
X"21",
X"21",
X"25",
X"27",
X"36",
X"2B",
X"2F",
X"36",
X"37",
X"3C",
X"25",
X"0E",
X"EC",
X"C9",
X"D0",
X"CA",
X"CC",
X"C4",
X"D0",
X"E5",
X"DE",
X"E4",
X"F7",
X"F7",
X"EB",
X"CD",
X"CF",
X"CD",
X"CD",
X"C9",
X"CD",
X"E5",
X"DB",
X"CB",
X"D3",
X"D9",
X"DC",
X"C5",
X"CD",
X"D1",
X"D9",
X"DD",
X"E4",
X"10",
X"26",
X"22",
X"29",
X"29",
X"2A",
X"13",
X"12",
X"15",
X"18",
X"1C",
X"0B",
X"1A",
X"27",
X"25",
X"2A",
X"24",
X"24",
X"07",
X"00",
X"FC",
X"F8",
X"0B",
X"0A",
X"18",
X"20",
X"15",
X"16",
X"0D",
X"0E",
X"F4",
X"E7",
X"E5",
X"C8",
X"C6",
X"C2",
X"D3",
X"E1",
X"D8",
X"DC",
X"D5",
X"DA",
X"C3",
X"BC",
X"DA",
X"DD",
X"E4",
X"E5",
X"F7",
X"0E",
X"0B",
X"13",
X"11",
X"1E",
X"06",
X"E2",
X"EE",
X"EF",
X"F7",
X"F6",
X"02",
X"1D",
X"1B",
X"22",
X"20",
X"36",
X"41",
X"26",
X"2B",
X"2B",
X"2C",
X"28",
X"29",
X"3B",
X"34",
X"31",
X"16",
X"06",
X"03",
X"E6",
X"E4",
X"E0",
X"DD",
X"DA",
X"DA",
X"EF",
X"F1",
X"01",
X"06",
X"00",
X"00",
X"E2",
X"DA",
X"DA",
X"D8",
X"D4",
X"D2",
X"E4",
X"D7",
X"D4",
X"DE",
X"E0",
X"EB",
X"D8",
X"D3",
X"DB",
X"E1",
X"E5",
X"ED",
X"12",
X"20",
X"1F",
X"24",
X"23",
X"2A",
X"1E",
X"15",
X"18",
X"1C",
X"16",
X"06",
X"16",
X"27",
X"27",
X"2C",
X"27",
X"28",
X"16",
X"04",
X"00",
X"07",
X"12",
X"08",
X"0D",
X"19",
X"12",
X"10",
X"0A",
X"08",
X"FE",
X"EA",
X"D7",
X"CA",
X"CC",
X"C8",
X"CC",
X"DD",
X"DC",
X"D9",
X"D7",
X"D6",
X"D0",
X"D1",
X"D8",
X"DB",
X"E2",
X"E6",
X"ED",
X"03",
X"09",
X"0C",
X"11",
X"10",
X"00",
X"F0",
X"F2",
X"F7",
X"FA",
X"FF",
X"01",
X"16",
X"20",
X"1E",
X"29",
X"3C",
X"3F",
X"2E",
X"27",
X"2D",
X"2B",
X"29",
X"23",
X"2C",
X"35",
X"20",
X"0D",
X"08",
X"07",
X"F6",
X"E6",
X"E7",
X"E3",
X"E1",
X"DD",
X"E4",
X"FE",
X"02",
X"00",
X"FA",
X"FA",
X"EC",
X"D8",
X"D9",
X"D5",
X"D5",
X"D1",
X"CA",
X"D4",
X"D9",
X"DF",
X"E3",
X"EA",
X"E8",
X"DA",
X"E0",
X"E5",
X"EB",
X"00",
X"0E",
X"22",
X"25",
X"27",
X"29",
X"2B",
X"2B",
X"18",
X"1B",
X"1B",
X"0B",
X"0B",
X"12",
X"27",
X"2D",
X"2D",
X"2C",
X"27",
X"22",
X"07",
X"04",
X"14",
X"0F",
X"0C",
X"07",
X"15",
X"16",
X"0F",
X"0D",
X"05",
X"06",
X"E9",
X"CD",
X"D0",
X"CB",
X"CC",
X"C8",
X"D7",
X"DF",
X"D8",
X"D9",
X"D2",
X"E0",
X"E0",
X"D4",
X"DF",
X"E1",
X"E8",
X"E9",
X"FC",
X"0C",
X"0B",
X"13",
X"03",
X"00",
X"FC",
X"F0",
X"F9",
X"FA",
X"00",
X"00",
X"0D",
X"20",
X"20",
X"36",
X"3E",
X"3F",
X"3A",
X"28",
X"2E",
X"2A",
X"2B",
X"23",
X"25",
X"30",
X"15",
X"0E",
X"09",
X"06",
X"00",
X"E9",
X"E8",
X"E2",
X"E2",
X"DC",
X"E2",
X"03",
X"01",
X"00",
X"FC",
X"F8",
X"F3",
X"DC",
X"D9",
X"D5",
X"D6",
X"CA",
X"B9",
X"D1",
X"D7",
X"DE",
X"E4",
X"E8",
X"EE",
X"DF",
X"DF",
X"E4",
X"F4",
X"07",
X"06",
X"1D",
X"26",
X"26",
X"2A",
X"2A",
X"2F",
X"1F",
X"1A",
X"11",
X"05",
X"0F",
X"0D",
X"20",
X"2D",
X"2D",
X"2C",
X"28",
X"24",
X"12",
X"11",
X"17",
X"0C",
X"0D",
X"03",
X"0D",
X"17",
X"10",
X"0C",
X"07",
X"03",
X"E5",
X"CD",
X"D0",
X"CA",
X"CE",
X"C6",
X"D0",
X"DD",
X"DC",
X"D6",
X"DE",
X"E9",
X"C5",
X"C8",
X"C9",
X"CC",
X"CE",
X"D0",
X"D1",
X"D4",
X"D6",
X"D7",
X"D9",
X"DB",
X"DD",
X"DE",
X"E0",
X"E1",
X"E2",
X"E3",
X"E5",
X"E6",
X"E7",
X"E8",
X"E9",
X"EA",
X"EB",
X"EC",
X"ED",
X"EE",
X"EF",
X"EF",
X"F0",
X"F0",
X"F1",
X"F2",
X"F3",
X"F3",
X"F4",
X"F4",
X"F5",
X"F5",
X"F6",
X"F5",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"0B",
X"09",
X"00",
X"FE",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FC",
X"FA",
X"FA",
X"FD",
X"00",
X"03",
X"07",
X"0A",
X"0D",
X"10",
X"14",
X"17",
X"1A",
X"1C",
X"1F",
X"21",
X"24",
X"26",
X"28",
X"2A",
X"2C",
X"2E",
X"30",
X"32",
X"33",
X"35",
X"36",
X"38",
X"39",
X"37",
X"33",
X"2C",
X"27",
X"21",
X"1C",
X"16",
X"12",
X"0D",
X"09",
X"04",
X"01",
X"FE",
X"FB",
X"F7",
X"F4",
X"F0",
X"ED",
X"EA",
X"E8",
X"E5",
X"E2",
X"DF",
X"DD",
X"DA",
X"D9",
X"D5",
X"D8",
X"D9",
X"DF",
X"E4",
X"E9",
X"EE",
X"F3",
X"F7",
X"FB",
X"FF",
X"01",
X"05",
X"08",
X"0C",
X"0F",
X"13",
X"16",
X"18",
X"1B",
X"1D",
X"20",
X"22",
X"24",
X"27",
X"2A",
X"2B",
X"2E",
X"2D",
X"2C",
X"26",
X"20",
X"1B",
X"16",
X"11",
X"0C",
X"08",
X"02",
X"00",
X"FD",
X"FA",
X"F6",
X"F6",
X"EE",
X"EF",
X"E6",
X"0C",
X"41",
X"33",
X"32",
X"27",
X"26",
X"17",
X"EE",
X"E9",
X"C4",
X"BA",
X"C2",
X"CC",
X"FC",
X"00",
X"05",
X"07",
X"0B",
X"0A",
X"EF",
X"10",
X"1D",
X"1A",
X"20",
X"1E",
X"4B",
X"53",
X"52",
X"51",
X"54",
X"4E",
X"03",
X"FA",
X"03",
X"01",
X"0A",
X"05",
X"2B",
X"35",
X"2C",
X"27",
X"2D",
X"4F",
X"26",
X"0C",
X"0E",
X"04",
X"06",
X"FC",
X"15",
X"24",
X"1F",
X"07",
X"E3",
X"ED",
X"CE",
X"B2",
X"B6",
X"B1",
X"B5",
X"AD",
X"C4",
X"DE",
X"F5",
X"0F",
X"02",
X"11",
X"00",
X"E5",
X"ED",
X"EF",
X"F8",
X"F6",
X"08",
X"0C",
X"FE",
X"09",
X"06",
X"10",
X"06",
X"E8",
X"EC",
X"F1",
X"F5",
X"FB",
X"2B",
X"5C",
X"59",
X"5C",
X"59",
X"5D",
X"53",
X"2B",
X"1E",
X"1F",
X"0F",
X"E7",
X"E3",
X"07",
X"09",
X"04",
X"00",
X"FF",
X"FA",
X"D4",
X"C1",
X"D5",
X"F2",
X"F0",
X"E9",
X"09",
X"14",
X"0A",
X"08",
X"03",
X"01",
X"E3",
X"B4",
X"9E",
X"A3",
X"AB",
X"AE",
X"D2",
X"F0",
X"EE",
X"F7",
X"F7",
X"FE",
X"03",
X"03",
X"08",
X"09",
X"10",
X"0B",
X"1F",
X"3D",
X"38",
X"3D",
X"3C",
X"24",
X"06",
X"F4",
X"FA",
X"FE",
X"01",
X"01",
X"0E",
X"2E",
X"20",
X"21",
X"3A",
X"40",
X"2A",
X"06",
X"02",
X"00",
X"FC",
X"F8",
X"FA",
X"1A",
X"0C",
X"E9",
X"E3",
X"E5",
X"DC",
X"B8",
X"B3",
X"B6",
X"B2",
X"B5",
X"B0",
X"E1",
X"00",
X"FE",
X"00",
X"02",
X"05",
X"EA",
X"E5",
X"EF",
X"EE",
X"F9",
X"E7",
X"F3",
X"03",
X"01",
X"0A",
X"0B",
X"11",
X"F8",
X"ED",
X"F8",
X"F5",
X"14",
X"27",
X"42",
X"57",
X"50",
X"54",
X"51",
X"55",
X"36",
X"1B",
X"1C",
X"F8",
X"EB",
X"E5",
X"F6",
X"0D",
X"00",
X"01",
X"FA",
X"FE",
X"E5",
X"C9",
X"ED",
X"EF",
X"ED",
X"E7",
X"F2",
X"0D",
X"02",
X"03",
X"FB",
X"FE",
X"E6",
X"A2",
X"A5",
X"A8",
X"AF",
X"B5",
X"C3",
X"EE",
X"ED",
X"F8",
X"F6",
X"09",
X"24",
X"03",
X"06",
X"0A",
X"0D",
X"11",
X"17",
X"3F",
X"3F",
X"44",
X"32",
X"18",
X"1E",
X"FE",
X"FD",
X"00",
X"02",
X"07",
X"05",
X"28",
X"27",
X"38",
X"49",
X"3A",
X"3B",
X"11",
X"02",
X"01",
X"FD",
X"F9",
X"ED",
X"03",
X"F5",
X"E1",
X"E6",
X"DD",
X"E1",
X"C5",
X"B4",
X"B7",
X"B4",
X"B7",
X"B3",
X"E4",
X"FB",
X"F2",
X"F9",
X"F9",
X"02",
X"F3",
X"E3",
X"EB",
X"EF",
X"F0",
X"D3",
X"E7",
X"04",
X"02",
X"0A",
X"09",
X"12",
X"06",
X"F4",
X"F8",
X"03",
X"24",
X"22",
X"2E",
X"4B",
X"4B",
X"4E",
X"4D",
X"4F",
X"41",
X"23",
X"0D",
X"F3",
X"F3",
X"ED",
X"EF",
X"07",
X"04",
X"00",
X"FE",
X"FD",
X"F3",
X"E7",
X"F3",
X"ED",
X"EA",
X"E5",
X"E6",
X"FF",
X"01",
X"FC",
X"FA",
X"F7",
X"DC",
X"AE",
X"AA",
X"AF",
X"B3",
X"BB",
X"C0",
X"E1",
X"F4",
X"F3",
X"FC",
X"17",
X"27",
X"0C",
X"03",
X"09",
X"0C",
X"0F",
X"10",
X"27",
X"3F",
X"36",
X"1E",
X"1A",
X"24",
X"10",
X"00",
X"06",
X"09",
X"0E",
X"0B",
X"16",
X"32",
X"44",
X"3F",
X"36",
X"33",
X"1F",
X"01",
X"00",
X"FC",
X"F8",
X"F6",
X"EE",
X"ED",
X"EB",
X"E9",
X"E5",
X"E4",
X"D9",
X"BB",
X"BA",
X"BA",
X"B7",
X"C8",
X"E2",
X"F8",
X"FB",
X"F9",
X"FF",
X"01",
X"02",
X"E9",
X"EB",
X"F3",
X"DE",
X"D5",
X"E0",
X"FC",
X"03",
X"04",
X"0B",
X"0C",
X"11",
X"FC",
X"FB",
X"16",
X"1F",
X"1F",
X"23",
X"3B",
X"47",
X"41",
X"47",
X"42",
X"44",
X"23",
X"FD",
X"FA",
X"F6",
X"F3",
X"EC",
X"FD",
X"08",
X"FF",
X"FF",
X"F6",
X"FF",
X"FF",
X"EB",
X"EC",
X"E7",
X"E7",
X"E1",
X"ED",
X"FF",
X"F4",
X"F8",
X"E4",
X"D2",
X"C4",
X"AF",
X"B7",
X"B9",
X"C3",
X"C5",
X"D7",
X"F4",
X"F1",
X"06",
X"19",
X"1B",
X"17",
X"01",
X"09",
X"0A",
X"0F",
X"10",
X"18",
X"36",
X"23",
X"19",
X"1E",
X"20",
X"20",
X"07",
X"0B",
X"0E",
X"11",
X"0F",
X"10",
X"3A",
X"3F",
X"35",
X"32",
X"29",
X"26",
X"06",
X"00",
X"FB",
X"F9",
X"F2",
X"D6",
X"E9",
X"F0",
X"E9",
X"E9",
X"E3",
X"E5",
X"C9",
X"C0",
X"BF",
X"C4",
X"DB",
X"D6",
X"E9",
X"F6",
X"F3",
X"FB",
X"FA",
X"02",
X"F2",
X"EC",
X"E7",
X"D5",
X"E0",
X"E0",
X"F6",
X"0A",
X"09",
X"11",
X"0F",
X"18",
X"09",
X"0A",
X"21",
X"1D",
X"25",
X"23",
X"31",
X"48",
X"45",
X"4A",
X"44",
X"47",
X"23",
X"FC",
X"FF",
X"F5",
X"F6",
X"EF",
X"F5",
X"06",
X"01",
X"00",
X"FD",
X"0E",
X"0C",
X"EE",
X"ED",
X"E9",
X"E7",
X"E3",
X"E5",
X"FA",
X"F9",
X"F2",
X"D7",
X"D2",
X"D1",
X"B5",
X"B6",
X"BA",
X"C3",
X"C8",
X"D0",
X"EC",
X"FF",
X"16",
X"1A",
X"1B",
X"20",
X"0A",
X"05",
X"0A",
X"0D",
X"10",
X"14",
X"21",
X"18",
X"1A",
X"1F",
X"1E",
X"25",
X"13",
X"09",
X"0F",
X"12",
X"10",
X"1A",
X"39",
X"3F",
X"36",
X"32",
X"29",
X"27",
X"12",
X"FE",
X"FD",
X"F9",
X"E5",
X"D0",
X"DF",
X"EF",
X"E9",
X"E9",
X"E5",
X"E5",
X"D8",
X"C0",
X"C1",
X"D4",
X"DC",
X"D4",
X"DD",
X"F3",
X"F2",
X"F8",
X"FD",
X"00",
X"00",
X"E9",
X"D7",
X"D8",
X"DF",
X"E1",
X"EC",
X"07",
X"0C",
X"0D",
X"14",
X"15",
X"1C",
X"1C",
X"1D",
X"20",
X"22",
X"23",
X"26",
X"41",
X"4A",
X"46",
X"4A",
X"3A",
X"20",
X"04",
X"FA",
X"F9",
X"F4",
X"F2",
X"ED",
X"FF",
X"06",
X"FC",
X"09",
X"15",
X"10",
X"FA",
X"E8",
X"EA",
X"E4",
X"E4",
X"DF",
X"EE",
X"FD",
X"E1",
X"D3",
X"D3",
X"D2",
X"C2",
X"B2",
X"BE",
X"C1",
X"CA",
X"CD",
X"DE",
X"04",
X"0B",
X"0E",
X"11",
X"16",
X"0F",
X"00",
X"09",
X"08",
X"0F",
X"0D",
X"05",
X"17",
X"1A",
X"1C",
X"20",
X"23",
X"21",
X"0E",
X"14",
X"13",
X"19",
X"28",
X"27",
X"36",
X"2F",
X"29",
X"23",
X"1E",
X"18",
X"FF",
X"FC",
X"F0",
X"DB",
X"DB",
X"D9",
X"EB",
X"EC",
X"E8",
X"E6",
X"E1",
X"E1",
X"C8",
X"CD",
X"DC",
X"D5",
X"D7",
X"D1",
X"E7",
X"EF",
X"F2",
X"F8",
X"F9",
X"00",
X"E4",
X"D5",
X"E0",
X"E2",
X"EB",
X"EB",
X"00",
X"0E",
X"0E",
X"13",
X"13",
X"2C",
X"26",
X"18",
X"21",
X"1E",
X"26",
X"22",
X"34",
X"43",
X"42",
X"41",
X"29",
X"23",
X"14",
X"FF",
X"00",
X"F9",
X"F9",
X"F0",
X"F8",
X"03",
X"01",
X"12",
X"0C",
X"0A",
X"00",
X"E9",
X"E9",
X"E3",
X"E4",
X"DD",
X"E3",
X"EB",
X"D7",
X"D7",
X"D4",
X"D2",
X"CF",
X"BC",
X"C1",
X"C7",
X"CF",
X"D2",
X"E4",
X"0B",
X"0E",
X"12",
X"15",
X"18",
X"1B",
X"09",
X"08",
X"0D",
X"11",
X"06",
X"FF",
X"18",
X"1F",
X"1F",
X"23",
X"23",
X"28",
X"18",
X"13",
X"18",
X"26",
X"2E",
X"21",
X"30",
X"31",
X"2A",
X"26",
X"1E",
X"1B",
X"08",
X"F9",
X"E6",
X"DC",
X"DF",
X"D7",
X"E4",
X"ED",
X"E8",
X"E7",
X"E3",
X"E1",
X"D7",
X"D9",
X"DC",
X"D6",
X"D8",
X"D1",
X"DE",
X"EE",
X"F2",
X"F7",
X"FC",
X"FB",
X"E5",
X"DA",
X"E1",
X"E4",
X"EB",
X"EC",
X"F8",
X"0C",
X"10",
X"11",
X"1F",
X"32",
X"2C",
X"1C",
X"1E",
X"20",
X"24",
X"24",
X"2B",
X"3E",
X"44",
X"34",
X"25",
X"24",
X"1C",
X"04",
X"FE",
X"FC",
X"F7",
X"F4",
X"F1",
X"00",
X"10",
X"12",
X"0C",
X"09",
X"04",
X"F1",
X"E6",
X"E7",
X"E1",
X"E1",
X"DB",
X"D8",
X"D9",
X"D6",
X"D5",
X"D2",
X"D2",
X"C6",
X"BE",
X"CB",
X"CC",
X"DA",
X"ED",
X"02",
X"10",
X"11",
X"14",
X"17",
X"1C",
X"13",
X"06",
X"10",
X"09",
X"FF",
X"00",
X"0D",
X"1F",
X"20",
X"23",
X"25",
X"28",
X"24",
X"11",
X"22",
X"2E",
X"2B",
X"23",
X"25",
X"31",
X"2A",
X"25",
X"1F",
X"1A",
X"12",
X"EE",
X"E0",
X"DF",
X"DD",
X"DA",
X"DA",
X"EC",
X"EA",
X"E7",
X"E4",
X"E1",
X"ED",
X"E3",
X"CD",
X"CB",
X"CD",
X"D0",
X"D1",
X"D4",
X"D6",
X"D8",
X"D9",
X"DB",
X"DC",
X"DE",
X"DF",
X"E1",
X"E2",
X"E4",
X"E5",
X"E6",
X"E8",
X"E9",
X"E9",
X"EB",
X"EB",
X"EC",
X"ED",
X"EE",
X"EF",
X"EF",
X"F0",
X"F1",
X"F1",
X"F2",
X"F3",
X"F3",
X"F4",
X"F4",
X"F5",
X"F6",
X"F6",
X"F6",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FE",
X"00",
X"1E",
X"1C",
X"02",
X"0F",
X"11",
X"0A",
X"03",
X"11",
X"11",
X"0E",
X"12",
X"11",
X"1B",
X"1B",
X"02",
X"00",
X"07",
X"00",
X"19",
X"F6",
X"03",
X"FE",
X"09",
X"00",
X"0F",
X"0E",
X"05",
X"04",
X"04",
X"02",
X"01",
X"02",
X"09",
X"0C",
X"12",
X"08",
X"04",
X"00",
X"04",
X"07",
X"19",
X"FE",
X"F3",
X"05",
X"F3",
X"00",
X"F5",
X"17",
X"F0",
X"00",
X"F9",
X"00",
X"00",
X"FF",
X"04",
X"04",
X"00",
X"00",
X"0B",
X"08",
X"00",
X"00",
X"03",
X"0A",
X"0D",
X"08",
X"F3",
X"F8",
X"F1",
X"02",
X"FB",
X"FF",
X"FF",
X"01",
X"13",
X"F8",
X"F9",
X"FF",
X"FA",
X"07",
X"05",
X"00",
X"FD",
X"FB",
X"FF",
X"FC",
X"03",
X"05",
X"0B",
X"0F",
X"03",
X"FB",
X"F7",
X"FF",
X"FD",
X"08",
X"FE",
X"FE",
X"05",
X"0D",
X"F5",
X"07",
X"09",
X"ED",
X"FF",
X"F6",
X"00",
X"FC",
X"09",
X"09",
X"FB",
X"02",
X"F9",
X"FB",
X"04",
X"00",
X"04",
X"03",
X"06",
X"0F",
X"01",
X"EE",
X"00",
X"F8",
X"06",
X"EE",
X"02",
X"FD",
X"FF",
X"FD",
X"01",
X"F2",
X"EA",
X"EE",
X"EC",
X"EF",
X"ED",
X"F2",
X"F0",
X"F2",
X"F1",
X"F3",
X"F2",
X"F4",
X"F3",
X"F4",
X"F5",
X"F6",
X"F6",
X"F6",
X"F7",
X"F8",
X"F6",
X"F9",
X"F8",
X"F9",
X"F9",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"03",
X"1D",
X"12",
X"18",
X"17",
X"0E",
X"16",
X"1A",
X"0B",
X"10",
X"0A",
X"09",
X"18",
X"1A",
X"FF",
X"0C",
X"0A",
X"01",
X"11",
X"0D",
X"00",
X"02",
X"10",
X"04",
X"00",
X"08",
X"0A",
X"0B",
X"02",
X"06",
X"08",
X"03",
X"04",
X"00",
X"F2",
X"E3",
X"F8",
X"F9",
X"F9",
X"F5",
X"01",
X"01",
X"0E",
X"08",
X"18",
X"1D",
X"1A",
X"12",
X"1C",
X"12",
X"1D",
X"23",
X"2A",
X"2B",
X"27",
X"3D",
X"35",
X"1E",
X"35",
X"30",
X"2A",
X"2B",
X"3F",
X"30",
X"21",
X"28",
X"1E",
X"2A",
X"14",
X"15",
X"1B",
X"0A",
X"FE",
X"09",
X"01",
X"01",
X"F3",
X"FA",
X"F7",
X"EC",
X"F4",
X"E2",
X"E2",
X"F0",
X"E5",
X"DF",
X"CE",
X"D6",
X"DB",
X"DA",
X"D4",
X"D2",
X"E2",
X"E7",
X"E6",
X"F3",
X"F7",
X"F9",
X"FB",
X"09",
X"00",
X"FA",
X"0A",
X"07",
X"14",
X"19",
X"1F",
X"1A",
X"13",
X"20",
X"28",
X"24",
X"12",
X"35",
X"28",
X"23",
X"31",
X"26",
X"32",
X"23",
X"27",
X"1F",
X"13",
X"0A",
X"14",
X"05",
X"FE",
X"FE",
X"F2",
X"F8",
X"F5",
X"01",
X"2F",
X"41",
X"40",
X"3F",
X"24",
X"28",
X"10",
X"EC",
X"FE",
X"D1",
X"BD",
X"B7",
X"C8",
X"F0",
X"02",
X"F2",
X"ED",
X"FE",
X"F2",
X"DB",
X"E4",
X"14",
X"0C",
X"1B",
X"19",
X"3E",
X"49",
X"51",
X"56",
X"46",
X"56",
X"03",
X"EF",
X"02",
X"FE",
X"01",
X"08",
X"37",
X"38",
X"38");
--//--------------------------------------
  begin

    if (RESET_N='0') then
      Q <= sqr_table(0);
    elsif(rising_edge(CLK)) then
      if (ENA='1') then
          Q <= sqr_table(to_integer(unsigned(ADDR)));
      end if;
    end if;
  end process;
end arch;