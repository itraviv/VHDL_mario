--------------------------------------
-- SinTable.vhd
-- Written by Saar Eliad and Itamar Raviv.
-- All rights reserved, Copyright 2017
--------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ThemeSoundTable is
port(
  CLK     : in std_logic;
  RESET_N : in std_logic;
  ENA     : in std_logic;
  ADDR    : in std_logic_vector(14 downto 0);
  Q       : out std_logic_vector(7 downto 0)
);
end ThemeSoundTable;

architecture arch of ThemeSoundTable is

type table_type is array(0 to 32767) of std_logic_vector(7 downto 0);
signal sqr_table : table_type;

begin

  SQRTableTC_proc: process(RESET_N, CLK)
    constant sqr_table : table_type := (

X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FE",
X"00",
X"FF",
X"01",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"02",
X"FD",
X"01",
X"FF",
X"00",
X"00",
X"02",
X"FA",
X"02",
X"FC",
X"03",
X"FB",
X"04",
X"FE",
X"07",
X"F8",
X"07",
X"F4",
X"10",
X"F9",
X"2C",
X"5A",
X"56",
X"4F",
X"4E",
X"4F",
X"37",
X"39",
X"2F",
X"38",
X"23",
X"2C",
X"1D",
X"3A",
X"0B",
X"0D",
X"09",
X"07",
X"06",
X"00",
X"01",
X"00",
X"00",
X"EA",
X"F7",
X"F2",
X"F7",
X"F2",
X"F7",
X"09",
X"14",
X"E9",
X"FC",
X"FC",
X"FE",
X"00",
X"09",
X"11",
X"0A",
X"1B",
X"0F",
X"2B",
X"11",
X"25",
X"19",
X"33",
X"22",
X"3F",
X"2E",
X"2C",
X"34",
X"27",
X"36",
X"39",
X"3B",
X"35",
X"34",
X"36",
X"24",
X"1A",
X"17",
X"0E",
X"14",
X"18",
X"1B",
X"F0",
X"F0",
X"F1",
X"E9",
X"00",
X"DB",
X"E2",
X"D8",
X"E8",
X"D7",
X"E1",
X"D6",
X"EA",
X"D5",
X"D0",
X"D2",
X"DF",
X"E0",
X"D8",
X"E7",
X"F9",
X"FB",
X"EF",
X"E7",
X"F5",
X"FF",
X"FB",
X"FF",
X"07",
X"11",
X"16",
X"15",
X"13",
X"35",
X"12",
X"10",
X"24",
X"1A",
X"2E",
X"1E",
X"2E",
X"26",
X"27",
X"2A",
X"35",
X"29",
X"24",
X"24",
X"1D",
X"1E",
X"10",
X"14",
X"0B",
X"04",
X"01",
X"0C",
X"F3",
X"F2",
X"EF",
X"EB",
X"E1",
X"F8",
X"E2",
X"E9",
X"D4",
X"09",
X"0F",
X"1C",
X"25",
X"17",
X"0E",
X"15",
X"1C",
X"14",
X"E7",
X"D4",
X"E2",
X"F4",
X"BD",
X"F1",
X"05",
X"14",
X"0F",
X"14",
X"1C",
X"24",
X"22",
X"1E",
X"31",
X"22",
X"34",
X"27",
X"65",
X"60",
X"6A",
X"62",
X"42",
X"34",
X"0C",
X"03",
X"00",
X"00",
X"FD",
X"ED",
X"20",
X"21",
X"08",
X"34",
X"35",
X"37",
X"10",
X"0E",
X"EC",
X"E2",
X"E4",
X"DC",
X"03",
X"0C",
X"EF",
X"CD",
X"E3",
X"DA",
X"B3",
X"99",
X"B1",
X"A9",
X"C1",
X"A5",
X"E2",
X"2D",
X"18",
X"23",
X"26",
X"2C",
X"1C",
X"09",
X"09",
X"FE",
X"05",
X"FE",
X"00",
X"1F",
X"18",
X"14",
X"1D",
X"36",
X"08",
X"E4",
X"01",
X"F1",
X"18",
X"26",
X"42",
X"5A",
X"60",
X"4B",
X"4D",
X"4A",
X"2B",
X"02",
X"0E",
X"F4",
X"CC",
X"C7",
X"D1",
X"FB",
X"F1",
X"F9",
X"EC",
X"EB",
X"E6",
X"B5",
X"DB",
X"EF",
X"DA",
X"E2",
X"E1",
X"05",
X"08",
X"10",
X"F8",
X"FA",
X"0D",
X"AB",
X"AB",
X"C5",
X"BA",
X"C8",
X"C1",
X"00",
X"16",
X"08",
X"0E",
X"1C",
X"3C",
X"25",
X"15",
X"1C",
X"0C",
X"2B",
X"13",
X"3C",
X"57",
X"54",
X"2C",
X"25",
X"20",
X"FC",
X"EE",
X"EE",
X"E2",
X"E8",
X"E9",
X"FF",
X"0F",
X"0B",
X"39",
X"25",
X"21",
X"0B",
X"E4",
X"F9",
X"F7",
X"F4",
X"CC",
X"E7",
X"E9",
X"CD",
X"E0",
X"C9",
X"D2",
X"C5",
X"B7",
X"9B",
X"A5",
X"AF",
X"B8",
X"E9",
X"07",
X"16",
X"1C",
X"18",
X"1D",
X"15",
X"0B",
X"0C",
X"FA",
X"0C",
X"F3",
X"F0",
X"12",
X"0B",
X"1F",
X"17",
X"2B",
X"20",
X"0A",
X"09",
X"F9",
X"23",
X"3B",
X"20",
X"52",
X"45",
X"54",
X"3F",
X"43",
X"31",
X"1B",
X"F8",
X"D8",
X"E1",
X"D8",
X"CB",
X"E8",
X"F0",
X"F4",
X"F6",
X"FF",
X"E0",
X"D4",
X"DB",
X"D8",
X"E0",
X"DF",
X"DD",
X"DC",
X"00",
X"F8",
X"FF",
X"00",
X"00",
X"D9",
X"B6",
X"AB",
X"C6",
X"CA",
X"C9",
X"D9",
X"04",
X"04",
X"14",
X"26",
X"34",
X"43",
X"0D",
X"0D",
X"1C",
X"16",
X"2E",
X"20",
X"44",
X"54",
X"1E",
X"1C",
X"28",
X"25",
X"03",
X"F4",
X"FF",
X"00",
X"EF",
X"F1",
X"11",
X"28",
X"37",
X"33",
X"2E",
X"11",
X"FE",
X"E8",
X"EB",
X"ED",
X"DD",
X"D7",
X"D6",
X"DD",
X"DA",
X"DC",
X"D7",
X"CE",
X"B9",
X"A2",
X"B9",
X"B4",
X"C7",
X"E4",
X"FA",
X"1B",
X"13",
X"05",
X"1B",
X"20",
X"04",
X"F8",
X"05",
X"F5",
X"EB",
X"FC",
X"FD",
X"14",
X"1B",
X"0A",
X"14",
X"18",
X"1D",
X"FD",
X"1A",
X"32",
X"3D",
X"25",
X"35",
X"4D",
X"3B",
X"3A",
X"27",
X"3A",
X"20",
X"EC",
X"DC",
X"DC",
X"E6",
X"DD",
X"D4",
X"00",
X"E0",
X"EC",
X"E9",
X"EB",
X"00",
X"DF",
X"E7",
X"E5",
X"D1",
X"D3",
X"DF",
X"F1",
X"00",
X"F9",
X"EB",
X"D8",
X"DF",
X"C7",
X"D3",
X"CA",
X"D0",
X"DF",
X"DB",
X"07",
X"19",
X"14",
X"29",
X"26",
X"2F",
X"22",
X"1D",
X"0B",
X"13",
X"1E",
X"20",
X"42",
X"2E",
X"22",
X"2D",
X"2D",
X"21",
X"16",
X"0D",
X"FC",
X"E5",
X"FC",
X"DB",
X"1F",
X"30",
X"16",
X"1B",
X"17",
X"16",
X"08",
X"EE",
X"E5",
X"EF",
X"E6",
X"C7",
X"D2",
X"DB",
X"D9",
X"E9",
X"DA",
X"E7",
X"CC",
X"B2",
X"B0",
X"B3",
X"E1",
X"ED",
X"FB",
X"0F",
X"14",
X"1C",
X"10",
X"27",
X"27",
X"EE",
X"FA",
X"DA",
X"E7",
X"EE",
X"FB",
X"0F",
X"0D",
X"16",
X"1B",
X"2C",
X"1F",
X"0A",
X"33",
X"28",
X"25",
X"3C",
X"31",
X"1E",
X"37",
X"1D",
X"2B",
X"19",
X"10",
X"EB",
X"D8",
X"DB",
X"D2",
X"D8",
X"D2",
X"EF",
X"E9",
X"F8",
X"ED",
X"00",
X"FC",
X"E5",
X"DB",
X"DF",
X"E3",
X"E8",
X"DA",
X"E0",
X"F3",
X"E0",
X"DC",
X"D7",
X"E6",
X"D8",
X"CD",
X"E0",
X"F0",
X"D1",
X"E0",
X"F1",
X"FD",
X"1D",
X"22",
X"2F",
X"27",
X"2B",
X"11",
X"2B",
X"07",
X"26",
X"1E",
X"27",
X"28",
X"26",
X"38",
X"35",
X"23",
X"1D",
X"FB",
X"03",
X"FA",
X"F7",
X"FF",
X"17",
X"3A",
X"1D",
X"16",
X"18",
X"12",
X"0C",
X"00",
X"D7",
X"E6",
X"DD",
X"C4",
X"C5",
X"D4",
X"DF",
X"D9",
X"E0",
X"D6",
X"DE",
X"C6",
X"AF",
X"C8",
X"E5",
X"E5",
X"E7",
X"05",
X"1C",
X"04",
X"13",
X"16",
X"18",
X"10",
X"EE",
X"EB",
X"E6",
X"F4",
X"FD",
X"09",
X"1B",
X"1C",
X"29",
X"31",
X"37",
X"21",
X"21",
X"25",
X"27",
X"36",
X"2B",
X"2F",
X"36",
X"37",
X"3C",
X"25",
X"0E",
X"EC",
X"C9",
X"D0",
X"CA",
X"CC",
X"C4",
X"D0",
X"E5",
X"DE",
X"E4",
X"F7",
X"F7",
X"EB",
X"CD",
X"CF",
X"CD",
X"CD",
X"C9",
X"CD",
X"E5",
X"DB",
X"CB",
X"D3",
X"D9",
X"DC",
X"C5",
X"CD",
X"D1",
X"D9",
X"DD",
X"E4",
X"10",
X"26",
X"22",
X"29",
X"29",
X"2A",
X"13",
X"12",
X"15",
X"18",
X"1C",
X"0B",
X"1A",
X"27",
X"25",
X"2A",
X"24",
X"24",
X"07",
X"00",
X"FC",
X"F8",
X"0B",
X"0A",
X"18",
X"20",
X"15",
X"16",
X"0D",
X"0E",
X"F4",
X"E7",
X"E5",
X"C8",
X"C6",
X"C2",
X"D3",
X"E1",
X"D8",
X"DC",
X"D5",
X"DA",
X"C3",
X"BC",
X"DA",
X"DD",
X"E4",
X"E5",
X"F7",
X"0E",
X"0B",
X"13",
X"11",
X"1E",
X"06",
X"E2",
X"EE",
X"EF",
X"F7",
X"F6",
X"02",
X"1D",
X"1B",
X"22",
X"20",
X"36",
X"41",
X"26",
X"2B",
X"2B",
X"2C",
X"28",
X"29",
X"3B",
X"34",
X"31",
X"16",
X"06",
X"03",
X"E6",
X"E4",
X"E0",
X"DD",
X"DA",
X"DA",
X"EF",
X"F1",
X"01",
X"06",
X"00",
X"00",
X"E2",
X"DA",
X"DA",
X"D8",
X"D4",
X"D2",
X"E4",
X"D7",
X"D4",
X"DE",
X"E0",
X"EB",
X"D8",
X"D3",
X"DB",
X"E1",
X"E5",
X"ED",
X"12",
X"20",
X"1F",
X"24",
X"23",
X"2A",
X"1E",
X"15",
X"18",
X"1C",
X"16",
X"06",
X"16",
X"27",
X"27",
X"2C",
X"27",
X"28",
X"16",
X"04",
X"00",
X"07",
X"12",
X"08",
X"0D",
X"19",
X"12",
X"10",
X"0A",
X"08",
X"FE",
X"EA",
X"D7",
X"CA",
X"CC",
X"C8",
X"CC",
X"DD",
X"DC",
X"D9",
X"D7",
X"D6",
X"D0",
X"D1",
X"D8",
X"DB",
X"E2",
X"E6",
X"ED",
X"03",
X"09",
X"0C",
X"11",
X"10",
X"00",
X"F0",
X"F2",
X"F7",
X"FA",
X"FF",
X"01",
X"16",
X"20",
X"1E",
X"29",
X"3C",
X"3F",
X"2E",
X"27",
X"2D",
X"2B",
X"29",
X"23",
X"2C",
X"35",
X"20",
X"0D",
X"08",
X"07",
X"F6",
X"E6",
X"E7",
X"E3",
X"E1",
X"DD",
X"E4",
X"FE",
X"02",
X"00",
X"FA",
X"FA",
X"EC",
X"D8",
X"D9",
X"D5",
X"D5",
X"D1",
X"CA",
X"D4",
X"D9",
X"DF",
X"E3",
X"EA",
X"E8",
X"DA",
X"E0",
X"E5",
X"EB",
X"00",
X"0E",
X"22",
X"25",
X"27",
X"29",
X"2B",
X"2B",
X"18",
X"1B",
X"1B",
X"0B",
X"0B",
X"12",
X"27",
X"2D",
X"2D",
X"2C",
X"27",
X"22",
X"07",
X"04",
X"14",
X"0F",
X"0C",
X"07",
X"15",
X"16",
X"0F",
X"0D",
X"05",
X"06",
X"E9",
X"CD",
X"D0",
X"CB",
X"CC",
X"C8",
X"D7",
X"DF",
X"D8",
X"D9",
X"D2",
X"E0",
X"E0",
X"D4",
X"DF",
X"E1",
X"E8",
X"E9",
X"FC",
X"0C",
X"0B",
X"13",
X"03",
X"00",
X"FC",
X"F0",
X"F9",
X"FA",
X"00",
X"00",
X"0D",
X"20",
X"20",
X"36",
X"3E",
X"3F",
X"3A",
X"28",
X"2E",
X"2A",
X"2B",
X"23",
X"25",
X"30",
X"15",
X"0E",
X"09",
X"06",
X"00",
X"E9",
X"E8",
X"E2",
X"E2",
X"DC",
X"E2",
X"03",
X"01",
X"00",
X"FC",
X"F8",
X"F3",
X"DC",
X"D9",
X"D5",
X"D6",
X"CA",
X"B9",
X"D1",
X"D7",
X"DE",
X"E4",
X"E8",
X"EE",
X"DF",
X"DF",
X"E4",
X"F4",
X"07",
X"06",
X"1D",
X"26",
X"26",
X"2A",
X"2A",
X"2F",
X"1F",
X"1A",
X"11",
X"05",
X"0F",
X"0D",
X"20",
X"2D",
X"2D",
X"2C",
X"28",
X"24",
X"12",
X"11",
X"17",
X"0C",
X"0D",
X"03",
X"0D",
X"17",
X"10",
X"0C",
X"07",
X"03",
X"E5",
X"CD",
X"D0",
X"CA",
X"CE",
X"C6",
X"D0",
X"DD",
X"DC",
X"D6",
X"DE",
X"E9",
X"C5",
X"C8",
X"C9",
X"CC",
X"CE",
X"D0",
X"D1",
X"D4",
X"D6",
X"D7",
X"D9",
X"DB",
X"DD",
X"DE",
X"E0",
X"E1",
X"E2",
X"E3",
X"E5",
X"E6",
X"E7",
X"E8",
X"E9",
X"EA",
X"EB",
X"EC",
X"ED",
X"EE",
X"EF",
X"EF",
X"F0",
X"F0",
X"F1",
X"F2",
X"F3",
X"F3",
X"F4",
X"F4",
X"F5",
X"F5",
X"F6",
X"F5",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"0B",
X"09",
X"00",
X"FE",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FC",
X"FA",
X"FA",
X"FD",
X"00",
X"03",
X"07",
X"0A",
X"0D",
X"10",
X"14",
X"17",
X"1A",
X"1C",
X"1F",
X"21",
X"24",
X"26",
X"28",
X"2A",
X"2C",
X"2E",
X"30",
X"32",
X"33",
X"35",
X"36",
X"38",
X"39",
X"37",
X"33",
X"2C",
X"27",
X"21",
X"1C",
X"16",
X"12",
X"0D",
X"09",
X"04",
X"01",
X"FE",
X"FB",
X"F7",
X"F4",
X"F0",
X"ED",
X"EA",
X"E8",
X"E5",
X"E2",
X"DF",
X"DD",
X"DA",
X"D9",
X"D5",
X"D8",
X"D9",
X"DF",
X"E4",
X"E9",
X"EE",
X"F3",
X"F7",
X"FB",
X"FF",
X"01",
X"05",
X"08",
X"0C",
X"0F",
X"13",
X"16",
X"18",
X"1B",
X"1D",
X"20",
X"22",
X"24",
X"27",
X"2A",
X"2B",
X"2E",
X"2D",
X"2C",
X"26",
X"20",
X"1B",
X"16",
X"11",
X"0C",
X"08",
X"02",
X"00",
X"FD",
X"FA",
X"F6",
X"F6",
X"EE",
X"EF",
X"E6",
X"0C",
X"41",
X"33",
X"32",
X"27",
X"26",
X"17",
X"EE",
X"E9",
X"C4",
X"BA",
X"C2",
X"CC",
X"FC",
X"00",
X"05",
X"07",
X"0B",
X"0A",
X"EF",
X"10",
X"1D",
X"1A",
X"20",
X"1E",
X"4B",
X"53",
X"52",
X"51",
X"54",
X"4E",
X"03",
X"FA",
X"03",
X"01",
X"0A",
X"05",
X"2B",
X"35",
X"2C",
X"27",
X"2D",
X"4F",
X"26",
X"0C",
X"0E",
X"04",
X"06",
X"FC",
X"15",
X"24",
X"1F",
X"07",
X"E3",
X"ED",
X"CE",
X"B2",
X"B6",
X"B1",
X"B5",
X"AD",
X"C4",
X"DE",
X"F5",
X"0F",
X"02",
X"11",
X"00",
X"E5",
X"ED",
X"EF",
X"F8",
X"F6",
X"08",
X"0C",
X"FE",
X"09",
X"06",
X"10",
X"06",
X"E8",
X"EC",
X"F1",
X"F5",
X"FB",
X"2B",
X"5C",
X"59",
X"5C",
X"59",
X"5D",
X"53",
X"2B",
X"1E",
X"1F",
X"0F",
X"E7",
X"E3",
X"07",
X"09",
X"04",
X"00",
X"FF",
X"FA",
X"D4",
X"C1",
X"D5",
X"F2",
X"F0",
X"E9",
X"09",
X"14",
X"0A",
X"08",
X"03",
X"01",
X"E3",
X"B4",
X"9E",
X"A3",
X"AB",
X"AE",
X"D2",
X"F0",
X"EE",
X"F7",
X"F7",
X"FE",
X"03",
X"03",
X"08",
X"09",
X"10",
X"0B",
X"1F",
X"3D",
X"38",
X"3D",
X"3C",
X"24",
X"06",
X"F4",
X"FA",
X"FE",
X"01",
X"01",
X"0E",
X"2E",
X"20",
X"21",
X"3A",
X"40",
X"2A",
X"06",
X"02",
X"00",
X"FC",
X"F8",
X"FA",
X"1A",
X"0C",
X"E9",
X"E3",
X"E5",
X"DC",
X"B8",
X"B3",
X"B6",
X"B2",
X"B5",
X"B0",
X"E1",
X"00",
X"FE",
X"00",
X"02",
X"05",
X"EA",
X"E5",
X"EF",
X"EE",
X"F9",
X"E7",
X"F3",
X"03",
X"01",
X"0A",
X"0B",
X"11",
X"F8",
X"ED",
X"F8",
X"F5",
X"14",
X"27",
X"42",
X"57",
X"50",
X"54",
X"51",
X"55",
X"36",
X"1B",
X"1C",
X"F8",
X"EB",
X"E5",
X"F6",
X"0D",
X"00",
X"01",
X"FA",
X"FE",
X"E5",
X"C9",
X"ED",
X"EF",
X"ED",
X"E7",
X"F2",
X"0D",
X"02",
X"03",
X"FB",
X"FE",
X"E6",
X"A2",
X"A5",
X"A8",
X"AF",
X"B5",
X"C3",
X"EE",
X"ED",
X"F8",
X"F6",
X"09",
X"24",
X"03",
X"06",
X"0A",
X"0D",
X"11",
X"17",
X"3F",
X"3F",
X"44",
X"32",
X"18",
X"1E",
X"FE",
X"FD",
X"00",
X"02",
X"07",
X"05",
X"28",
X"27",
X"38",
X"49",
X"3A",
X"3B",
X"11",
X"02",
X"01",
X"FD",
X"F9",
X"ED",
X"03",
X"F5",
X"E1",
X"E6",
X"DD",
X"E1",
X"C5",
X"B4",
X"B7",
X"B4",
X"B7",
X"B3",
X"E4",
X"FB",
X"F2",
X"F9",
X"F9",
X"02",
X"F3",
X"E3",
X"EB",
X"EF",
X"F0",
X"D3",
X"E7",
X"04",
X"02",
X"0A",
X"09",
X"12",
X"06",
X"F4",
X"F8",
X"03",
X"24",
X"22",
X"2E",
X"4B",
X"4B",
X"4E",
X"4D",
X"4F",
X"41",
X"23",
X"0D",
X"F3",
X"F3",
X"ED",
X"EF",
X"07",
X"04",
X"00",
X"FE",
X"FD",
X"F3",
X"E7",
X"F3",
X"ED",
X"EA",
X"E5",
X"E6",
X"FF",
X"01",
X"FC",
X"FA",
X"F7",
X"DC",
X"AE",
X"AA",
X"AF",
X"B3",
X"BB",
X"C0",
X"E1",
X"F4",
X"F3",
X"FC",
X"17",
X"27",
X"0C",
X"03",
X"09",
X"0C",
X"0F",
X"10",
X"27",
X"3F",
X"36",
X"1E",
X"1A",
X"24",
X"10",
X"00",
X"06",
X"09",
X"0E",
X"0B",
X"16",
X"32",
X"44",
X"3F",
X"36",
X"33",
X"1F",
X"01",
X"00",
X"FC",
X"F8",
X"F6",
X"EE",
X"ED",
X"EB",
X"E9",
X"E5",
X"E4",
X"D9",
X"BB",
X"BA",
X"BA",
X"B7",
X"C8",
X"E2",
X"F8",
X"FB",
X"F9",
X"FF",
X"01",
X"02",
X"E9",
X"EB",
X"F3",
X"DE",
X"D5",
X"E0",
X"FC",
X"03",
X"04",
X"0B",
X"0C",
X"11",
X"FC",
X"FB",
X"16",
X"1F",
X"1F",
X"23",
X"3B",
X"47",
X"41",
X"47",
X"42",
X"44",
X"23",
X"FD",
X"FA",
X"F6",
X"F3",
X"EC",
X"FD",
X"08",
X"FF",
X"FF",
X"F6",
X"FF",
X"FF",
X"EB",
X"EC",
X"E7",
X"E7",
X"E1",
X"ED",
X"FF",
X"F4",
X"F8",
X"E4",
X"D2",
X"C4",
X"AF",
X"B7",
X"B9",
X"C3",
X"C5",
X"D7",
X"F4",
X"F1",
X"06",
X"19",
X"1B",
X"17",
X"01",
X"09",
X"0A",
X"0F",
X"10",
X"18",
X"36",
X"23",
X"19",
X"1E",
X"20",
X"20",
X"07",
X"0B",
X"0E",
X"11",
X"0F",
X"10",
X"3A",
X"3F",
X"35",
X"32",
X"29",
X"26",
X"06",
X"00",
X"FB",
X"F9",
X"F2",
X"D6",
X"E9",
X"F0",
X"E9",
X"E9",
X"E3",
X"E5",
X"C9",
X"C0",
X"BF",
X"C4",
X"DB",
X"D6",
X"E9",
X"F6",
X"F3",
X"FB",
X"FA",
X"02",
X"F2",
X"EC",
X"E7",
X"D5",
X"E0",
X"E0",
X"F6",
X"0A",
X"09",
X"11",
X"0F",
X"18",
X"09",
X"0A",
X"21",
X"1D",
X"25",
X"23",
X"31",
X"48",
X"45",
X"4A",
X"44",
X"47",
X"23",
X"FC",
X"FF",
X"F5",
X"F6",
X"EF",
X"F5",
X"06",
X"01",
X"00",
X"FD",
X"0E",
X"0C",
X"EE",
X"ED",
X"E9",
X"E7",
X"E3",
X"E5",
X"FA",
X"F9",
X"F2",
X"D7",
X"D2",
X"D1",
X"B5",
X"B6",
X"BA",
X"C3",
X"C8",
X"D0",
X"EC",
X"FF",
X"16",
X"1A",
X"1B",
X"20",
X"0A",
X"05",
X"0A",
X"0D",
X"10",
X"14",
X"21",
X"18",
X"1A",
X"1F",
X"1E",
X"25",
X"13",
X"09",
X"0F",
X"12",
X"10",
X"1A",
X"39",
X"3F",
X"36",
X"32",
X"29",
X"27",
X"12",
X"FE",
X"FD",
X"F9",
X"E5",
X"D0",
X"DF",
X"EF",
X"E9",
X"E9",
X"E5",
X"E5",
X"D8",
X"C0",
X"C1",
X"D4",
X"DC",
X"D4",
X"DD",
X"F3",
X"F2",
X"F8",
X"FD",
X"00",
X"00",
X"E9",
X"D7",
X"D8",
X"DF",
X"E1",
X"EC",
X"07",
X"0C",
X"0D",
X"14",
X"15",
X"1C",
X"1C",
X"1D",
X"20",
X"22",
X"23",
X"26",
X"41",
X"4A",
X"46",
X"4A",
X"3A",
X"20",
X"04",
X"FA",
X"F9",
X"F4",
X"F2",
X"ED",
X"FF",
X"06",
X"FC",
X"09",
X"15",
X"10",
X"FA",
X"E8",
X"EA",
X"E4",
X"E4",
X"DF",
X"EE",
X"FD",
X"E1",
X"D3",
X"D3",
X"D2",
X"C2",
X"B2",
X"BE",
X"C1",
X"CA",
X"CD",
X"DE",
X"04",
X"0B",
X"0E",
X"11",
X"16",
X"0F",
X"00",
X"09",
X"08",
X"0F",
X"0D",
X"05",
X"17",
X"1A",
X"1C",
X"20",
X"23",
X"21",
X"0E",
X"14",
X"13",
X"19",
X"28",
X"27",
X"36",
X"2F",
X"29",
X"23",
X"1E",
X"18",
X"FF",
X"FC",
X"F0",
X"DB",
X"DB",
X"D9",
X"EB",
X"EC",
X"E8",
X"E6",
X"E1",
X"E1",
X"C8",
X"CD",
X"DC",
X"D5",
X"D7",
X"D1",
X"E7",
X"EF",
X"F2",
X"F8",
X"F9",
X"00",
X"E4",
X"D5",
X"E0",
X"E2",
X"EB",
X"EB",
X"00",
X"0E",
X"0E",
X"13",
X"13",
X"2C",
X"26",
X"18",
X"21",
X"1E",
X"26",
X"22",
X"34",
X"43",
X"42",
X"41",
X"29",
X"23",
X"14",
X"FF",
X"00",
X"F9",
X"F9",
X"F0",
X"F8",
X"03",
X"01",
X"12",
X"0C",
X"0A",
X"00",
X"E9",
X"E9",
X"E3",
X"E4",
X"DD",
X"E3",
X"EB",
X"D7",
X"D7",
X"D4",
X"D2",
X"CF",
X"BC",
X"C1",
X"C7",
X"CF",
X"D2",
X"E4",
X"0B",
X"0E",
X"12",
X"15",
X"18",
X"1B",
X"09",
X"08",
X"0D",
X"11",
X"06",
X"FF",
X"18",
X"1F",
X"1F",
X"23",
X"23",
X"28",
X"18",
X"13",
X"18",
X"26",
X"2E",
X"21",
X"30",
X"31",
X"2A",
X"26",
X"1E",
X"1B",
X"08",
X"F9",
X"E6",
X"DC",
X"DF",
X"D7",
X"E4",
X"ED",
X"E8",
X"E7",
X"E3",
X"E1",
X"D7",
X"D9",
X"DC",
X"D6",
X"D8",
X"D1",
X"DE",
X"EE",
X"F2",
X"F7",
X"FC",
X"FB",
X"E5",
X"DA",
X"E1",
X"E4",
X"EB",
X"EC",
X"F8",
X"0C",
X"10",
X"11",
X"1F",
X"32",
X"2C",
X"1C",
X"1E",
X"20",
X"24",
X"24",
X"2B",
X"3E",
X"44",
X"34",
X"25",
X"24",
X"1C",
X"04",
X"FE",
X"FC",
X"F7",
X"F4",
X"F1",
X"00",
X"10",
X"12",
X"0C",
X"09",
X"04",
X"F1",
X"E6",
X"E7",
X"E1",
X"E1",
X"DB",
X"D8",
X"D9",
X"D6",
X"D5",
X"D2",
X"D2",
X"C6",
X"BE",
X"CB",
X"CC",
X"DA",
X"ED",
X"02",
X"10",
X"11",
X"14",
X"17",
X"1C",
X"13",
X"06",
X"10",
X"09",
X"FF",
X"00",
X"0D",
X"1F",
X"20",
X"23",
X"25",
X"28",
X"24",
X"11",
X"22",
X"2E",
X"2B",
X"23",
X"25",
X"31",
X"2A",
X"25",
X"1F",
X"1A",
X"12",
X"EE",
X"E0",
X"DF",
X"DD",
X"DA",
X"DA",
X"EC",
X"EA",
X"E7",
X"E4",
X"E1",
X"ED",
X"E3",
X"CD",
X"CB",
X"CD",
X"D0",
X"D1",
X"D4",
X"D6",
X"D8",
X"D9",
X"DB",
X"DC",
X"DE",
X"DF",
X"E1",
X"E2",
X"E4",
X"E5",
X"E6",
X"E8",
X"E9",
X"E9",
X"EB",
X"EB",
X"EC",
X"ED",
X"EE",
X"EF",
X"EF",
X"F0",
X"F1",
X"F1",
X"F2",
X"F3",
X"F3",
X"F4",
X"F4",
X"F5",
X"F6",
X"F6",
X"F6",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FE",
X"00",
X"1E",
X"1C",
X"02",
X"0F",
X"11",
X"0A",
X"03",
X"11",
X"11",
X"0E",
X"12",
X"11",
X"1B",
X"1B",
X"02",
X"00",
X"07",
X"00",
X"19",
X"F6",
X"03",
X"FE",
X"09",
X"00",
X"0F",
X"0E",
X"05",
X"04",
X"04",
X"02",
X"01",
X"02",
X"09",
X"0C",
X"12",
X"08",
X"04",
X"00",
X"04",
X"07",
X"19",
X"FE",
X"F3",
X"05",
X"F3",
X"00",
X"F5",
X"17",
X"F0",
X"00",
X"F9",
X"00",
X"00",
X"FF",
X"04",
X"04",
X"00",
X"00",
X"0B",
X"08",
X"00",
X"00",
X"03",
X"0A",
X"0D",
X"08",
X"F3",
X"F8",
X"F1",
X"02",
X"FB",
X"FF",
X"FF",
X"01",
X"13",
X"F8",
X"F9",
X"FF",
X"FA",
X"07",
X"05",
X"00",
X"FD",
X"FB",
X"FF",
X"FC",
X"03",
X"05",
X"0B",
X"0F",
X"03",
X"FB",
X"F7",
X"FF",
X"FD",
X"08",
X"FE",
X"FE",
X"05",
X"0D",
X"F5",
X"07",
X"09",
X"ED",
X"FF",
X"F6",
X"00",
X"FC",
X"09",
X"09",
X"FB",
X"02",
X"F9",
X"FB",
X"04",
X"00",
X"04",
X"03",
X"06",
X"0F",
X"01",
X"EE",
X"00",
X"F8",
X"06",
X"EE",
X"02",
X"FD",
X"FF",
X"FD",
X"01",
X"F2",
X"EA",
X"EE",
X"EC",
X"EF",
X"ED",
X"F2",
X"F0",
X"F2",
X"F1",
X"F3",
X"F2",
X"F4",
X"F3",
X"F4",
X"F5",
X"F6",
X"F6",
X"F6",
X"F7",
X"F8",
X"F6",
X"F9",
X"F8",
X"F9",
X"F9",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"03",
X"1D",
X"12",
X"18",
X"17",
X"0E",
X"16",
X"1A",
X"0B",
X"10",
X"0A",
X"09",
X"18",
X"1A",
X"FF",
X"0C",
X"0A",
X"01",
X"11",
X"0D",
X"00",
X"02",
X"10",
X"04",
X"00",
X"08",
X"0A",
X"0B",
X"02",
X"06",
X"08",
X"03",
X"04",
X"00",
X"F2",
X"E3",
X"F8",
X"F9",
X"F9",
X"F5",
X"01",
X"01",
X"0E",
X"08",
X"18",
X"1D",
X"1A",
X"12",
X"1C",
X"12",
X"1D",
X"23",
X"2A",
X"2B",
X"27",
X"3D",
X"35",
X"1E",
X"35",
X"30",
X"2A",
X"2B",
X"3F",
X"30",
X"21",
X"28",
X"1E",
X"2A",
X"14",
X"15",
X"1B",
X"0A",
X"FE",
X"09",
X"01",
X"01",
X"F3",
X"FA",
X"F7",
X"EC",
X"F4",
X"E2",
X"E2",
X"F0",
X"E5",
X"DF",
X"CE",
X"D6",
X"DB",
X"DA",
X"D4",
X"D2",
X"E2",
X"E7",
X"E6",
X"F3",
X"F7",
X"F9",
X"FB",
X"09",
X"00",
X"FA",
X"0A",
X"07",
X"14",
X"19",
X"1F",
X"1A",
X"13",
X"20",
X"28",
X"24",
X"12",
X"35",
X"28",
X"23",
X"31",
X"26",
X"32",
X"23",
X"27",
X"1F",
X"13",
X"0A",
X"14",
X"05",
X"FE",
X"FE",
X"F2",
X"F8",
X"F5",
X"01",
X"2F",
X"41",
X"40",
X"3F",
X"24",
X"28",
X"10",
X"EC",
X"FE",
X"D1",
X"BD",
X"B7",
X"C8",
X"F0",
X"02",
X"F2",
X"ED",
X"FE",
X"F2",
X"DB",
X"E4",
X"14",
X"0C",
X"1B",
X"19",
X"3E",
X"49",
X"51",
X"56",
X"46",
X"56",
X"03",
X"EF",
X"02",
X"FE",
X"01",
X"08",
X"37",
X"38",
X"27",
X"39",
X"28",
X"41",
X"37",
X"18",
X"17",
X"0C",
X"17",
X"12",
X"2A",
X"21",
X"28",
X"1F",
X"F4",
X"E8",
X"D9",
X"B1",
X"B7",
X"B9",
X"B7",
X"C4",
X"D1",
X"D8",
X"EC",
X"03",
X"06",
X"0D",
X"F0",
X"CD",
X"E5",
X"E4",
X"EC",
X"EA",
X"FF",
X"16",
X"FD",
X"02",
X"08",
X"02",
X"F8",
X"E5",
X"E8",
X"EF",
X"F4",
X"EC",
X"0C",
X"5F",
X"49",
X"5B",
X"5C",
X"62",
X"4E",
X"1C",
X"20",
X"25",
X"32",
X"05",
X"DA",
X"15",
X"12",
X"12",
X"00",
X"04",
X"0B",
X"D2",
X"C9",
X"CE",
X"F4",
X"0B",
X"DC",
X"0A",
X"16",
X"06",
X"11",
X"F9",
X"0E",
X"D5",
X"D0",
X"9F",
X"A9",
X"A4",
X"A4",
X"C7",
X"D9",
X"E8",
X"ED",
X"EB",
X"F8",
X"E3",
X"FE",
X"0F",
X"01",
X"00",
X"00",
X"14",
X"40",
X"3F",
X"39",
X"32",
X"2E",
X"FD",
X"E8",
X"08",
X"FD",
X"EE",
X"ED",
X"00",
X"24",
X"2A",
X"28",
X"28",
X"46",
X"3E",
X"0D",
X"0E",
X"0D",
X"13",
X"17",
X"04",
X"12",
X"25",
X"ED",
X"DE",
X"DD",
X"E0",
X"AA",
X"B9",
X"AD",
X"C8",
X"B8",
X"B7",
X"D7",
X"FB",
X"01",
X"00",
X"04",
X"00",
X"E5",
X"D4",
X"D6",
X"E6",
X"EA",
X"E9",
X"F7",
X"FF",
X"0A",
X"00",
X"01",
X"0E",
X"EB",
X"E5",
X"04",
X"F0",
X"E7",
X"1E",
X"34",
X"50",
X"45",
X"46",
X"41",
X"59",
X"3E",
X"1A",
X"2E",
X"1D",
X"01",
X"F5",
X"10",
X"15",
X"16",
X"14",
X"09",
X"07",
X"FF",
X"C3",
X"DB",
X"01",
X"FA",
X"DE",
X"F7",
X"05",
X"0A",
X"03",
X"FF",
X"FC",
X"00",
X"C5",
X"93",
X"AD",
X"9D",
X"AD",
X"B3",
X"EC",
X"EE",
X"DB",
X"EA",
X"E8",
X"07",
X"00",
X"01",
X"08",
X"07",
X"06",
X"11",
X"2E",
X"34",
X"3D",
X"47",
X"21",
X"0F",
X"FF",
X"FD",
X"F2",
X"08",
X"0A",
X"FC",
X"26",
X"2F",
X"2E",
X"57",
X"4E",
X"42",
X"1D",
X"14",
X"03",
X"04",
X"02",
X"FF",
X"14",
X"09",
X"F0",
X"EE",
X"E5",
X"F3",
X"CE",
X"C0",
X"BA",
X"C0",
X"CC",
X"C4",
X"D9",
X"F6",
X"EE",
X"F1",
X"F5",
X"FC",
X"E3",
X"CD",
X"E5",
X"E0",
X"EE",
X"D3",
X"D5",
X"FE",
X"FD",
X"FD",
X"07",
X"16",
X"FC",
X"E5",
X"F8",
X"F1",
X"0C",
X"32",
X"2F",
X"38",
X"43",
X"35",
X"4A",
X"40",
X"49",
X"22",
X"1D",
X"0C",
X"FC",
X"F7",
X"04",
X"23",
X"0B",
X"11",
X"01",
X"07",
X"FD",
X"E8",
X"FE",
X"F7",
X"F3",
X"F7",
X"E3",
X"0B",
X"0D",
X"F5",
X"00",
X"F7",
X"F3",
X"BB",
X"BA",
X"BA",
X"A6",
X"9C",
X"AC",
X"D8",
X"DA",
X"DB",
X"E6",
X"FC",
X"23",
X"FE",
X"F8",
X"10",
X"0D",
X"F5",
X"02",
X"0C",
X"3E",
X"2F",
X"1C",
X"07",
X"17",
X"08",
X"F5",
X"04",
X"02",
X"17",
X"FA",
X"27",
X"2C",
X"4C",
X"55",
X"38",
X"50",
X"35",
X"0A",
X"09",
X"06",
X"03",
X"F8",
X"13",
X"05",
X"EE",
X"FD",
X"EE",
X"F1",
X"EA",
X"D5",
X"AB",
X"C5",
X"C0",
X"B4",
X"D8",
X"FE",
X"F4",
X"F1",
X"F4",
X"F2",
X"F7",
X"E1",
X"E4",
X"E6",
X"E0",
X"C7",
X"D9",
X"F0",
X"0D",
X"00",
X"F4",
X"04",
X"F8",
X"F5",
X"ED",
X"14",
X"18",
X"00",
X"23",
X"24",
X"3B",
X"31",
X"4B",
X"42",
X"3A",
X"28",
X"13",
X"02",
X"02",
X"01",
X"FD",
X"11",
X"20",
X"0A",
X"0F",
X"06",
X"FA",
X"00",
X"FE",
X"03",
X"E9",
X"F3",
X"F0",
X"EF",
X"FB",
X"F9",
X"03",
X"F0",
X"DA",
X"D1",
X"BE",
X"A8",
X"B3",
X"AD",
X"C1",
X"CA",
X"DB",
X"EF",
X"E0",
X"08",
X"12",
X"06",
X"00",
X"05",
X"04",
X"16",
X"FE",
X"0B",
X"36",
X"21",
X"1F",
X"11",
X"21",
X"13",
X"00",
X"0A",
X"11",
X"15",
X"14",
X"1D",
X"3A",
X"48",
X"4F",
X"49",
X"3C",
X"20",
X"0E",
X"07",
X"09",
X"FB",
X"02",
X"EC",
X"F4",
X"FD",
X"F7",
X"F6",
X"F0",
X"DA",
X"CB",
X"C7",
X"CD",
X"C5",
X"BE",
X"DD",
X"E2",
X"FC",
X"E9",
X"F2",
X"01",
X"EC",
X"D7",
X"D0",
X"D9",
X"D8",
X"C8",
X"DC",
X"E5",
X"0E",
X"F8",
X"06",
X"00",
X"14",
X"02",
X"01",
X"23",
X"15",
X"22",
X"1B",
X"21",
X"49",
X"4A",
X"45",
X"40",
X"44",
X"3E",
X"0E",
X"F6",
X"F1",
X"EE",
X"E8",
X"F0",
X"02",
X"FA",
X"F9",
X"F3",
X"FE",
X"05",
X"E8",
X"EB",
X"E5",
X"E4",
X"DE",
X"E3",
X"F6",
X"F0",
X"F1",
X"DF",
X"CB",
X"CC",
X"AF",
X"AE",
X"AD",
X"B0",
X"B1",
X"BB",
X"DA",
X"E4",
X"F8",
X"09",
X"07",
X"10",
X"FB",
X"FA",
X"FE",
X"01",
X"05",
X"06",
X"20",
X"16",
X"0D",
X"16",
X"13",
X"1C",
X"06",
X"01",
X"06",
X"0A",
X"0D",
X"11",
X"3C",
X"4D",
X"40",
X"3E",
X"34",
X"33",
X"19",
X"06",
X"04",
X"00",
X"FA",
X"DC",
X"E8",
X"F9",
X"EF",
X"F1",
X"E9",
X"EC",
X"DC",
X"C6",
X"C5",
X"CC",
X"E1",
X"DB",
X"E2",
X"F7",
X"EF",
X"EF",
X"ED",
X"F4",
X"ED",
X"DF",
X"D6",
X"C9",
X"D3",
X"D5",
X"E1",
X"00",
X"01",
X"06",
X"08",
X"0E",
X"0A",
X"07",
X"18",
X"17",
X"1C",
X"1D",
X"21",
X"3D",
X"43",
X"41",
X"44",
X"45",
X"30",
X"0B",
X"08",
X"03",
X"00",
X"FE",
X"FB",
X"0A",
X"10",
X"07",
X"07",
X"19",
X"1C",
X"00",
X"F3",
X"F1",
X"ED",
X"EB",
X"E7",
X"F8",
X"02",
X"F5",
X"DE",
X"D7",
X"DA",
X"C3",
X"B5",
X"B6",
X"B7",
X"BA",
X"BF",
X"D0",
X"ED",
X"00",
X"03",
X"05",
X"0C",
X"02",
X"F9",
X"FF",
X"02",
X"05",
X"09",
X"0A",
X"0F",
X"12",
X"15",
X"18",
X"1D",
X"17",
X"08",
X"0C",
X"10",
X"11",
X"22",
X"35",
X"43",
X"3F",
X"37",
X"31",
X"2B",
X"21",
X"09",
X"04",
X"00",
X"ED",
X"E1",
X"E4",
X"F4",
X"F3",
X"EE",
X"ED",
X"E9",
X"E6",
X"CE",
X"CB",
X"DE",
X"DF",
X"DB",
X"D9",
X"EA",
X"EE",
X"E7",
X"EB",
X"EA",
X"F4",
X"DF",
X"CB",
X"D4",
X"DA",
X"DF",
X"E2",
X"F8",
X"05",
X"03",
X"0B",
X"0A",
X"19",
X"1C",
X"12",
X"18",
X"1A",
X"1F",
X"1E",
X"2E",
X"3F",
X"3A",
X"40",
X"32",
X"2A",
X"1F",
X"0D",
X"0C",
X"05",
X"03",
X"FE",
X"03",
X"11",
X"06",
X"13",
X"17",
X"13",
X"06",
X"F2",
X"F3",
X"EE",
X"ED",
X"E7",
X"EA",
X"FB",
X"E4",
X"DB",
X"DA",
X"D8",
X"D2",
X"BC",
X"BC",
X"BC",
X"C1",
X"C5",
X"D0",
X"FC",
X"03",
X"05",
X"0A",
X"0C",
X"0F",
X"FF",
X"00",
X"03",
X"08",
X"08",
X"FA",
X"0E",
X"16",
X"17",
X"1C",
X"1C",
X"21",
X"0F",
X"0F",
X"11",
X"19",
X"30",
X"2D",
X"3D",
X"41",
X"37",
X"34",
X"2A",
X"29",
X"10",
X"05",
X"FA",
X"E6",
X"E9",
X"E1",
X"EE",
X"F6",
X"EF",
X"F0",
X"E9",
X"EB",
X"D8",
X"D6",
X"E4",
X"DB",
X"DD",
X"D6",
X"E2",
X"ED",
X"E8",
X"EB",
X"EA",
X"F4",
X"DD",
X"C9",
X"D6",
X"D7",
X"E0",
X"E1",
X"F0",
X"04",
X"05",
X"0A",
X"0D",
X"25",
X"25",
X"12",
X"19",
X"19",
X"1E",
X"1E",
X"26",
X"3A",
X"3D",
X"3B",
X"28",
X"2A",
X"27",
X"11",
X"0B",
X"06",
X"03",
X"00",
X"FE",
X"0A",
X"10",
X"1C",
X"17",
X"12",
X"0E",
X"F8",
X"F1",
X"EE",
X"EB",
X"E7",
X"E6",
X"EB",
X"DF",
X"DD",
X"DB",
X"D8",
X"D8",
X"C4",
X"BA",
X"BE",
X"BF",
X"C5",
X"D7",
X"F9",
X"03",
X"05",
X"0A",
X"0B",
X"12",
X"06",
X"FF",
X"04",
X"07",
X"FD",
X"F5",
X"07",
X"18",
X"18",
X"1B",
X"1D",
X"22",
X"1A",
X"0C",
X"13",
X"26",
X"30",
X"2C",
X"34",
X"41",
X"39",
X"33",
X"2C",
X"28",
X"1C",
X"01",
X"EE",
X"E8",
X"E7",
X"E1",
X"E6",
X"F5",
X"F2",
X"EE",
X"ED",
X"E6",
X"EC",
X"E0",
X"D0",
X"D7",
X"D6",
X"DA",
X"DA",
X"DD",
X"DD",
X"DF",
X"E0",
X"E2",
X"E2",
X"E4",
X"E5",
X"E7",
X"E8",
X"E9",
X"EA",
X"EB",
X"EB",
X"EC",
X"ED",
X"EE",
X"EF",
X"F0",
X"F0",
X"F1",
X"F2",
X"F2",
X"F4",
X"F4",
X"F4",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F7",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FE",
X"00",
X"FF",
X"00",
X"FE",
X"00",
X"FC",
X"07",
X"15",
X"14",
X"10",
X"02",
X"16",
X"0B",
X"0D",
X"0C",
X"1B",
X"21",
X"0E",
X"00",
X"09",
X"02",
X"0C",
X"0F",
X"0F",
X"00",
X"08",
X"0E",
X"14",
X"0C",
X"01",
X"13",
X"0B",
X"00",
X"09",
X"13",
X"FA",
X"FF",
X"F5",
X"ED",
X"F9",
X"F1",
X"F8",
X"E5",
X"ED",
X"F2",
X"ED",
X"ED",
X"00",
X"00",
X"F4",
X"04",
X"FA",
X"FF",
X"02",
X"13",
X"15",
X"15",
X"1E",
X"29",
X"27",
X"17",
X"1F",
X"14",
X"29",
X"1E",
X"34",
X"26",
X"2D",
X"3B",
X"2E",
X"2D",
X"3F",
X"36",
X"23",
X"19",
X"11",
X"1D",
X"12",
X"11",
X"06",
X"0C",
X"14",
X"FD",
X"FF",
X"F8",
X"F4",
X"FE",
X"02",
X"DE",
X"DF",
X"E5",
X"CF",
X"EA",
X"D9",
X"D2",
X"CE",
X"DA",
X"D0",
X"D9",
X"CB",
X"E0",
X"EA",
X"ED",
X"E7",
X"F0",
X"F7",
X"01",
X"F8",
X"06",
X"0B",
X"F8",
X"09",
X"04",
X"1B",
X"12",
X"14",
X"24",
X"1E",
X"16",
X"23",
X"26",
X"32",
X"2A",
X"19",
X"2D",
X"25",
X"3C",
X"1C",
X"22",
X"1D",
X"16",
X"0D",
X"18",
X"1C",
X"04",
X"FD",
X"E8",
X"02",
X"13",
X"08",
X"08",
X"00",
X"0D",
X"29",
X"1D",
X"1C",
X"12",
X"13",
X"EA",
X"DD",
X"BF",
X"A9",
X"AD",
X"B0",
X"B7",
X"BA",
X"C1",
X"CA",
X"FE",
X"26",
X"30",
X"2E",
X"34",
X"30",
X"38",
X"25",
X"09",
X"10",
X"13",
X"10",
X"EE",
X"F2",
X"F4",
X"17",
X"2C",
X"27",
X"2E",
X"2B",
X"31",
X"2F",
X"39",
X"2F",
X"28",
X"23",
X"21",
X"16",
X"15",
X"0A",
X"1F",
X"36",
X"2F",
X"15",
X"F2",
X"F7",
X"EC",
X"F1",
X"C4",
X"B8",
X"B9",
X"B8",
X"BB",
X"B4",
X"D0",
X"EA",
X"0A",
X"08",
X"03",
X"00",
X"01",
X"01",
X"0B",
X"F8",
X"DF",
X"C9",
X"BB",
X"CA",
X"CA",
X"D7",
X"D5",
X"01",
X"0D",
X"11",
X"14",
X"19",
X"40",
X"4D",
X"41",
X"1C",
X"20",
X"21",
X"24",
X"27",
X"29",
X"29",
X"3B",
X"2F",
X"22",
X"22",
X"18",
X"18",
X"0E",
X"10",
X"E2",
X"D8",
X"D3",
X"E0",
X"00",
X"FD",
X"F7",
X"FF",
X"1F",
X"19",
X"15",
X"10",
X"0B",
X"09",
X"F5",
X"B6",
X"A0",
X"A4",
X"A3",
X"A4",
X"A7",
X"AD",
X"B2",
X"E2",
X"EC",
X"09",
X"27",
X"21",
X"1D",
X"1D",
X"17",
X"F8",
X"00",
X"01",
X"06",
X"0A",
X"F5",
X"E5",
X"06",
X"1C",
X"1D",
X"20",
X"22",
X"24",
X"25",
X"26",
X"08",
X"23",
X"2C",
X"24",
X"21",
X"1A",
X"15",
X"1A",
X"38",
X"2B",
X"2C",
X"1C",
X"FB",
X"F0",
X"F4",
X"D2",
X"BF",
X"C0",
X"C0",
X"BE",
X"BF",
X"B9",
X"C7",
X"06",
X"05",
X"01",
X"FF",
X"FB",
X"F8",
X"FB",
X"F0",
X"D3",
X"E3",
X"D1",
X"BE",
X"C6",
X"CE",
X"CF",
X"F3",
X"06",
X"06",
X"0A",
X"0F",
X"0E",
X"2B",
X"40",
X"18",
X"1C",
X"1B",
X"21",
X"21",
X"25",
X"24",
X"36",
X"59",
X"35",
X"25",
X"26",
X"1D",
X"1B",
X"17",
X"F8",
X"E2",
X"E5",
X"DF",
X"E0",
X"FD",
X"00",
X"FE",
X"20",
X"18",
X"17",
X"0D",
X"0D",
X"04",
X"08",
X"EC",
X"AB",
X"AC",
X"AB",
X"AD",
X"AC",
X"AC",
X"AE",
X"CE",
X"E6",
X"E1",
X"F5",
X"16",
X"18",
X"1C",
X"19",
X"F9",
X"FF",
X"00",
X"06",
X"04",
X"12",
X"FD",
X"FB",
X"1B",
X"18",
X"1F",
X"1D",
X"22",
X"24",
X"28",
X"0C",
X"FF",
X"1E",
X"34",
X"2D",
X"2A",
X"1F",
X"23",
X"36",
X"2F",
X"29",
X"1F",
X"1F",
X"00",
X"F4",
X"E3",
X"C6",
X"CC",
X"C6",
X"C9",
X"C5",
X"C4",
X"C2",
X"DE",
X"00",
X"00",
X"FA",
X"F9",
X"F2",
X"F4",
X"E8",
X"D0",
X"D2",
X"D8",
X"DB",
X"C3",
X"C8",
X"CB",
X"E6",
X"00",
X"FE",
X"04",
X"01",
X"0C",
X"0B",
X"19",
X"19",
X"15",
X"19",
X"1B",
X"1D",
X"22",
X"20",
X"2F",
X"49",
X"4B",
X"40",
X"26",
X"2A",
X"24",
X"23",
X"08",
X"F1",
X"F3",
X"EB",
X"EE",
X"E4",
X"F8",
X"04",
X"1A",
X"1D",
X"14",
X"12",
X"0D",
X"08",
X"08",
X"F8",
X"DC",
X"C4",
X"B2",
X"B8",
X"B2",
X"B6",
X"AF",
X"C7",
X"D8",
X"D7",
X"E0",
X"E3",
X"04",
X"10",
X"0E",
X"F8",
X"F5",
X"FD",
X"FF",
X"02",
X"05",
X"07",
X"13",
X"14",
X"10",
X"18",
X"16",
X"1F",
X"1C",
X"25",
X"0C",
X"03",
X"06",
X"12",
X"32",
X"2F",
X"2D",
X"2A",
X"40",
X"3F",
X"36",
X"32",
X"2A",
X"28",
X"17",
X"ED",
X"D3",
X"D3",
X"D0",
X"D1",
X"CC",
X"CD",
X"C7",
X"E1",
X"E8",
X"F6",
X"06",
X"FE",
X"FF",
X"F9",
X"F3",
X"D1",
X"CE",
X"D1",
X"D2",
X"D7",
X"C9",
X"C0",
X"D8",
X"EF",
X"F2",
X"F7",
X"FA",
X"00",
X"00",
X"06",
X"F6",
X"04",
X"13",
X"11",
X"18",
X"17",
X"1D",
X"20",
X"3E",
X"3E",
X"42",
X"3E",
X"29",
X"25",
X"29",
X"16",
X"00",
X"00",
X"FB",
X"F8",
X"F3",
X"EF",
X"F1",
X"1A",
X"1D",
X"16",
X"13",
X"0D",
X"0B",
X"04",
X"00",
X"E1",
X"E3",
X"D3",
X"BD",
X"BE",
X"BD",
X"B9",
X"C7",
X"D8",
X"D1",
X"D6",
X"D7",
X"DC",
X"F0",
X"06",
X"F0",
X"F0",
X"F5",
X"F8",
X"FC",
X"00",
X"02",
X"09",
X"28",
X"14",
X"0C",
X"13",
X"14",
X"17",
X"1C",
X"10",
X"01",
X"0A",
X"09",
X"10",
X"27",
X"34",
X"2D",
X"46",
X"43",
X"3D",
X"36",
X"32",
X"29",
X"27",
X"17",
X"E4",
X"E0",
X"DE",
X"DC",
X"D9",
X"D8",
X"D3",
X"E1",
X"F1",
X"E6",
X"EE",
X"00",
X"FE",
X"F8",
X"F7",
X"D8",
X"D4",
X"D0",
X"D2",
X"D1",
X"DA",
X"D2",
X"CA",
X"EB",
X"EB",
X"F4",
X"F5",
X"FC",
X"FD",
X"03",
X"F7",
X"E9",
X"01",
X"13",
X"14",
X"17",
X"1A",
X"1D",
X"38",
X"3D",
X"3F",
X"3E",
X"43",
X"2E",
X"25",
X"23",
X"07",
X"0C",
X"02",
X"03",
X"FC",
X"FD",
X"F5",
X"03",
X"24",
X"23",
X"1D",
X"18",
X"12",
X"0E",
X"08",
X"ED",
X"E6",
X"E5",
X"E0",
X"C4",
X"C1",
X"BF",
X"C6",
X"DD",
X"D5",
X"D9",
X"D1",
X"D7",
X"D3",
X"E5",
X"ED",
X"E5",
X"ED",
X"F0",
X"F5",
X"F9",
X"FD",
X"02",
X"1D",
X"25",
X"1B",
X"09",
X"0F",
X"0F",
X"15",
X"0E",
X"FD",
X"05",
X"02",
X"0B",
X"08",
X"20",
X"2F",
X"44",
X"4F",
X"48",
X"44",
X"3B",
X"35",
X"2F",
X"27",
X"0A",
X"F3",
X"E1",
X"E4",
X"DD",
X"DF",
X"D7",
X"E3",
X"F4",
X"ED",
X"ED",
X"E7",
X"FE",
X"FF",
X"FC",
X"E3",
X"D6",
X"D8",
X"D2",
X"D3",
X"D1",
X"D4",
X"D8",
X"E0",
X"E0",
X"EA",
X"EB",
X"F3",
X"F3",
X"FD",
X"F1",
X"E4",
X"EA",
X"F4",
X"11",
X"11",
X"17",
X"17",
X"31",
X"3C",
X"39",
X"3F",
X"3E",
X"41",
X"37",
X"1F",
X"0A",
X"0D",
X"0A",
X"0B",
X"04",
X"04",
X"FB",
X"08",
X"12",
X"19",
X"29",
X"1D",
X"1D",
X"14",
X"13",
X"F6",
X"EB",
X"EC",
X"E6",
X"E7",
X"D0",
X"C0",
X"C7",
X"DE",
X"D8",
X"D4",
X"D2",
X"D2",
X"CD",
X"D3",
X"C5",
X"D0",
X"E0",
X"E1",
X"EA",
X"EB",
X"F3",
X"F4",
X"0C",
X"14",
X"18",
X"19",
X"08",
X"08",
X"0E",
X"0B",
X"FD",
X"00",
X"03",
X"07",
X"0A",
X"0D",
X"12",
X"37",
X"46",
X"45",
X"45",
X"40",
X"3C",
X"33",
X"30",
X"13",
X"0D",
X"00",
X"EE",
X"EC",
X"E8",
X"E3",
X"E8",
X"F9",
X"F4",
X"F0",
X"EC",
X"E8",
X"F0",
X"FF",
X"E8",
X"DB",
X"DB",
X"D8",
X"D7",
X"D3",
X"D3",
X"D1",
X"EA",
X"E2",
X"DC",
X"E3",
X"E7",
X"ED",
X"F2",
X"EF",
X"E1",
X"E8",
X"EC",
X"F2",
X"04",
X"12",
X"0F",
X"24",
X"2F",
X"2F",
X"32",
X"32",
X"35",
X"37",
X"35",
X"10",
X"0C",
X"11",
X"14",
X"14",
X"12",
X"0B",
X"0F",
X"1C",
X"13",
X"14",
X"20",
X"1F",
X"17",
X"15",
X"00",
X"F4",
X"F3",
X"EF",
X"EC",
X"EB",
X"E0",
X"CD",
X"E1",
X"E0",
X"DD",
X"DA",
X"D8",
X"D5",
X"D5",
X"CB",
X"B9",
X"CB",
X"E0",
X"E3",
X"E8",
X"EE",
X"F0",
X"03",
X"11",
X"12",
X"15",
X"18",
X"0D",
X"04",
X"0A",
X"F9",
X"FD",
X"00",
X"04",
X"05",
X"0B",
X"0A",
X"19",
X"3C",
X"44",
X"43",
X"44",
X"43",
X"3F",
X"3A",
X"23",
X"15",
X"13",
X"0C",
X"F7",
X"EF",
X"EE",
X"EC",
X"FE",
X"FA",
X"F9",
X"F2",
X"F3",
X"EB",
X"EF",
X"F4",
X"E3",
X"E2",
X"DE",
X"DE",
X"DA",
X"D9",
X"D6",
X"E4",
X"ED",
X"E4",
X"D6",
X"DD",
X"E2",
X"E7",
X"E9",
X"D9",
X"DF",
X"E2",
X"EB",
X"EC",
X"FE",
X"0C",
X"19",
X"2C",
X"2A",
X"2E",
X"2E",
X"31",
X"32",
X"34",
X"24",
X"12",
X"0A",
X"10",
X"11",
X"16",
X"14",
X"17",
X"24",
X"1E",
X"1B",
X"13",
X"22",
X"23",
X"1E",
X"0D",
X"FB",
X"FC",
X"F5",
X"F5",
X"EF",
X"EF",
X"E8",
X"E7",
X"E3",
X"E2",
X"DE",
X"DE",
X"D9",
X"DA",
X"D0",
X"BD",
X"BB",
X"C1",
X"D8",
X"DE",
X"E4",
X"E8",
X"FA",
X"0A",
X"08",
X"0F",
X"0F",
X"16",
X"10",
X"03",
X"F4",
X"F5",
X"F9",
X"FE",
X"00",
X"05",
X"05",
X"12",
X"24",
X"30",
X"42",
X"40",
X"43",
X"42",
X"44",
X"31",
X"20",
X"1E",
X"15",
X"15",
X"02",
X"F3",
X"F2",
X"00",
X"00",
X"FD",
X"FA",
X"F7",
X"F2",
X"F2",
X"E8",
X"D9",
X"DF",
X"DD",
X"E1",
X"E0",
X"E3",
X"E3",
X"E6",
X"E6",
X"E8",
X"E8",
X"EA",
X"EB",
X"EC",
X"ED",
X"EE",
X"EE",
X"EF",
X"F0",
X"F1",
X"F1",
X"F2",
X"F2",
X"F3",
X"F3",
X"F4",
X"F4",
X"F5",
X"F6",
X"F6",
X"F6",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"01",
X"00",
X"00",
X"FE",
X"08",
X"14",
X"0A",
X"18",
X"0F",
X"16",
X"0E",
X"0D",
X"0C",
X"14",
X"1D",
X"0B",
X"11",
X"09",
X"04",
X"07",
X"0F",
X"0A",
X"0B",
X"13",
X"18",
X"03",
X"05",
X"00",
X"FD",
X"08",
X"01",
X"03",
X"02",
X"14",
X"09",
X"F8",
X"F3",
X"F0",
X"F7",
X"00",
X"E1",
X"E1",
X"E2",
X"E0",
X"E6",
X"E6",
X"E9",
X"E8",
X"E0",
X"EE",
X"EA",
X"FD",
X"00",
X"02",
X"07",
X"01",
X"0D",
X"0C",
X"1A",
X"18",
X"0C",
X"1B",
X"20",
X"24",
X"17",
X"27",
X"29",
X"21",
X"36",
X"24",
X"2E",
X"38",
X"2B",
X"35",
X"32",
X"1B",
X"28",
X"1D",
X"0D",
X"12",
X"10",
X"11",
X"02",
X"00",
X"02",
X"ED",
X"EB",
X"F5",
X"F0",
X"F0",
X"E6",
X"EF",
X"F3",
X"D3",
X"E0",
X"D8",
X"D5",
X"D3",
X"E0",
X"DD",
X"C4",
X"E4",
X"D3",
X"DD",
X"EC",
X"E1",
X"F0",
X"F5",
X"F7",
X"01",
X"08",
X"FD",
X"17",
X"06",
X"08",
X"10",
X"13",
X"1E",
X"1F",
X"2B",
X"27",
X"16",
X"19",
X"1F",
X"27",
X"40",
X"1F",
X"27",
X"23",
X"21",
X"1C",
X"1B",
X"21",
X"10",
X"0A",
X"23",
X"41",
X"60",
X"4B",
X"49",
X"49",
X"3B",
X"2A",
X"0A",
X"F2",
X"E6",
X"C2",
X"C3",
X"D8",
X"F8",
X"F3",
X"DD",
X"E7",
X"E0",
X"E2",
X"AA",
X"D5",
X"FF",
X"FC",
X"FB",
X"0E",
X"2D",
X"34",
X"35",
X"32",
X"38",
X"2F",
X"F5",
X"E4",
X"E4",
X"F5",
X"EF",
X"F4",
X"34",
X"24",
X"23",
X"34",
X"36",
X"4F",
X"2E",
X"2A",
X"32",
X"2C",
X"31",
X"31",
X"4D",
X"55",
X"45",
X"30",
X"10",
X"0B",
X"CD",
X"CC",
X"D3",
X"C5",
X"D5",
X"D2",
X"F1",
X"F1",
X"EE",
X"22",
X"11",
X"08",
X"F3",
X"D2",
X"DC",
X"E0",
X"DC",
X"CF",
X"F3",
X"EF",
X"DC",
X"DE",
X"E1",
X"EF",
X"D2",
X"CB",
X"D2",
X"C0",
X"E6",
X"D0",
X"15",
X"45",
X"33",
X"48",
X"47",
X"43",
X"2F",
X"1E",
X"28",
X"19",
X"27",
X"00",
X"00",
X"36",
X"26",
X"2F",
X"2B",
X"2A",
X"1A",
X"F3",
X"E6",
X"DF",
X"07",
X"1E",
X"09",
X"2E",
X"2B",
X"25",
X"24",
X"28",
X"12",
X"E9",
X"D9",
X"AD",
X"B3",
X"B7",
X"C0",
X"DA",
X"D9",
X"E9",
X"D3",
X"CC",
X"D7",
X"AF",
X"D2",
X"E3",
X"E9",
X"E7",
X"E2",
X"18",
X"17",
X"18",
X"22",
X"28",
X"14",
X"EB",
X"E7",
X"DD",
X"DE",
X"F0",
X"E0",
X"18",
X"25",
X"18",
X"1E",
X"3A",
X"5A",
X"47",
X"1E",
X"23",
X"21",
X"1A",
X"10",
X"32",
X"44",
X"29",
X"1E",
X"FF",
X"18",
X"E8",
X"C6",
X"DD",
X"D0",
X"BF",
X"C8",
X"DD",
X"EB",
X"FE",
X"10",
X"01",
X"0B",
X"F0",
X"D0",
X"DC",
X"DD",
X"D1",
X"CD",
X"E0",
X"DC",
X"CC",
X"E8",
X"EA",
X"E6",
X"DF",
X"C2",
X"D2",
X"E1",
X"E3",
X"DD",
X"15",
X"37",
X"36",
X"43",
X"31",
X"3F",
X"43",
X"28",
X"0E",
X"29",
X"15",
X"EB",
X"01",
X"24",
X"2B",
X"2A",
X"39",
X"32",
X"1F",
X"EF",
X"E8",
X"FA",
X"14",
X"0C",
X"01",
X"22",
X"29",
X"21",
X"21",
X"2C",
X"05",
X"F2",
X"C9",
X"A6",
X"B4",
X"AE",
X"B3",
X"C4",
X"EF",
X"D9",
X"DB",
X"D0",
X"CD",
X"DE",
X"D3",
X"E9",
X"E2",
X"F0",
X"FA",
X"0E",
X"12",
X"24",
X"21",
X"0E",
X"0D",
X"ED",
X"D3",
X"DE",
X"E9",
X"F6",
X"F2",
X"FB",
X"35",
X"30",
X"20",
X"49",
X"52",
X"45",
X"31",
X"2D",
X"2D",
X"24",
X"21",
X"22",
X"3C",
X"25",
X"12",
X"08",
X"FB",
X"F4",
X"DB",
X"D0",
X"D1",
X"D8",
X"C8",
X"C9",
X"FD",
X"0D",
X"08",
X"00",
X"03",
X"04",
X"DB",
X"CF",
X"DC",
X"D6",
X"CF",
X"C0",
X"CB",
X"CF",
X"D8",
X"E1",
X"E7",
X"F7",
X"DD",
X"D5",
X"E0",
X"DC",
X"FA",
X"0E",
X"1C",
X"39",
X"33",
X"37",
X"3A",
X"39",
X"24",
X"1F",
X"20",
X"02",
X"FF",
X"00",
X"16",
X"3A",
X"30",
X"1D",
X"27",
X"22",
X"09",
X"F3",
X"08",
X"12",
X"0E",
X"15",
X"01",
X"22",
X"17",
X"0A",
X"10",
X"0E",
X"F2",
X"B9",
X"D3",
X"C3",
X"B2",
X"B9",
X"B0",
X"EA",
X"D8",
X"D4",
X"C8",
X"DD",
X"FA",
X"DD",
X"DF",
X"E3",
X"ED",
X"FE",
X"FA",
X"09",
X"15",
X"14",
X"07",
X"05",
X"0F",
X"E8",
X"E2",
X"FB",
X"F5",
X"EE",
X"F6",
X"18",
X"2B",
X"35",
X"4F",
X"55",
X"50",
X"33",
X"1F",
X"29",
X"2F",
X"1F",
X"17",
X"23",
X"1A",
X"1B",
X"0A",
X"F6",
X"0B",
X"E0",
X"DF",
X"D7",
X"D0",
X"C8",
X"D4",
X"08",
X"10",
X"05",
X"0B",
X"01",
X"06",
X"ED",
X"DE",
X"D4",
X"D7",
X"C1",
X"AE",
X"C0",
X"E4",
X"CF",
X"E8",
X"DF",
X"EB",
X"E8",
X"DC",
X"D7",
X"F4",
X"11",
X"07",
X"09",
X"28",
X"1B",
X"27",
X"2B",
X"35",
X"28",
X"1D",
X"16",
X"16",
X"F3",
X"FA",
X"01",
X"17",
X"2A",
X"14",
X"28",
X"09",
X"1A",
X"00",
X"1E",
X"FF",
X"0E",
X"FF",
X"06",
X"06",
X"23",
X"14",
X"03",
X"04",
X"ED",
X"D7",
X"CA",
X"C6",
X"C5",
X"C4",
X"C9",
X"E4",
X"EB",
X"D0",
X"D4",
X"ED",
X"F5",
X"FA",
X"C7",
X"D5",
X"E0",
X"DD",
X"F2",
X"F6",
X"20",
X"0C",
X"05",
X"F7",
X"04",
X"FA",
X"EF",
X"F7",
X"F8",
X"0E",
X"0A",
X"0C",
X"2C",
X"46",
X"4C",
X"41",
X"4D",
X"4E",
X"21",
X"34",
X"20",
X"1D",
X"2C",
X"08",
X"0C",
X"15",
X"0A",
X"17",
X"03",
X"EF",
X"DF",
X"CB",
X"DE",
X"D2",
X"E6",
X"F0",
X"08",
X"08",
X"03",
X"01",
X"EC",
X"F9",
X"DF",
X"DD",
X"CF",
X"B5",
X"B9",
X"C2",
X"DF",
X"E6",
X"ED",
X"E9",
X"ED",
X"F5",
X"E6",
X"F3",
X"FE",
X"06",
X"09",
X"01",
X"23",
X"3D",
X"35",
X"28",
X"31",
X"3F",
X"1C",
X"E9",
X"EF",
X"F2",
X"F8",
X"FC",
X"0D",
X"21",
X"19",
X"19",
X"0A",
X"1D",
X"15",
X"02",
X"01",
X"FC",
X"FA",
X"F4",
X"FD",
X"0E",
X"02",
X"06",
X"ED",
X"DF",
X"D5",
X"BA",
X"BC",
X"BA",
X"BC",
X"B9",
X"C1",
X"D7",
X"D1",
X"E8",
X"EC",
X"ED",
X"EB",
X"D7",
X"DF",
X"E2",
X"E9",
X"EC",
X"F5",
X"11",
X"FD",
X"FC",
X"00",
X"04",
X"04",
X"F0",
X"F3",
X"F7",
X"FD",
X"00",
X"06",
X"3A",
X"43",
X"41",
X"45",
X"41",
X"45",
X"2D",
X"26",
X"23",
X"20",
X"14",
X"F7",
X"0C",
X"0D",
X"06",
X"06",
X"00",
X"00",
X"E6",
X"DB",
X"D8",
X"E2",
X"F5",
X"EA",
X"FE",
X"05",
X"FF",
X"FD",
X"F6",
X"F9",
X"E0",
X"D1",
X"C2",
X"AE",
X"B8",
X"B4",
X"CC",
X"E4",
X"E6",
X"EE",
X"EF",
X"F9",
X"EE",
X"F3",
X"05",
X"00",
X"09",
X"08",
X"17",
X"2E",
X"2D",
X"31",
X"32",
X"35",
X"17",
X"FE",
X"05",
X"05",
X"0B",
X"0B",
X"18",
X"2F",
X"2D",
X"27",
X"25",
X"39",
X"31",
X"11",
X"0C",
X"07",
X"04",
X"00",
X"00",
X"11",
X"13",
X"05",
X"EC",
X"EA",
X"E6",
X"CB",
X"C5",
X"C5",
X"C4",
X"C2",
X"C1",
X"D0",
X"DF",
X"EA",
X"E7",
X"E8",
X"EC",
X"E0",
X"DC",
X"E6",
X"E8",
X"EE",
X"F2",
X"FA",
X"FA",
X"FE",
X"01",
X"03",
X"09",
X"00",
X"F7",
X"00",
X"00",
X"05",
X"16",
X"30",
X"3C",
X"3B",
X"3D",
X"3D",
X"40",
X"37",
X"24",
X"27",
X"1C",
X"08",
X"FD",
X"04",
X"0F",
X"08",
X"05",
X"00",
X"FF",
X"F5",
X"DE",
X"E2",
X"F1",
X"F2",
X"EB",
X"EF",
X"FE",
X"FA",
X"F5",
X"F3",
X"EF",
X"EB",
X"CC",
X"BA",
X"B8",
X"BC",
X"BE",
X"C8",
X"E1",
X"E9",
X"EC",
X"F2",
X"F3",
X"00",
X"00",
X"00",
X"04",
X"07",
X"0C",
X"0F",
X"24",
X"2C",
X"2A",
X"31",
X"23",
X"1A",
X"0C",
X"08",
X"0F",
X"0F",
X"14",
X"15",
X"28",
X"2F",
X"25",
X"32",
X"33",
X"2D",
X"19",
X"08",
X"09",
X"01",
X"00",
X"F9",
X"03",
X"0B",
X"F4",
X"ED",
X"EB",
X"E9",
X"DA",
X"C8",
X"CB",
X"C6",
X"C9",
X"C2",
X"D0",
X"F1",
X"ED",
X"EB",
X"EB",
X"F0",
X"ED",
X"DF",
X"E8",
X"E9",
X"F2",
X"ED",
X"E7",
X"FE",
X"00",
X"04",
X"07",
X"0B",
X"0B",
X"FB",
X"00",
X"00",
X"0F",
X"21",
X"26",
X"3D",
X"3E",
X"3E",
X"40",
X"41",
X"41",
X"29",
X"27",
X"15",
X"02",
X"01",
X"FE",
X"0C",
X"0C",
X"06",
X"02",
X"FF",
X"FE",
X"E5",
X"ED",
X"F7",
X"EF",
X"EF",
X"E9",
X"F8",
X"FB",
X"F5",
X"F4",
X"EF",
X"EE",
X"C7",
X"B7",
X"BB",
X"B9",
X"C0",
X"C2",
X"DA",
X"E8",
X"EB",
X"F1",
X"F7",
X"10",
X"07",
X"FF",
X"06",
X"06",
X"0B",
X"0A",
X"1D",
X"2C",
X"2D",
X"2A",
X"19",
X"1F",
X"16",
X"08",
X"10",
X"11",
X"16",
X"15",
X"20",
X"2E",
X"30",
X"3B",
X"32",
X"2F",
X"22",
X"0A",
X"07",
X"02",
X"00",
X"FA",
X"FF",
X"00",
X"EF",
X"EF",
X"E9",
X"E9",
X"E2",
X"CD",
X"CA",
X"C8",
X"C8",
X"C4",
X"D4",
X"F0",
X"EC",
X"EB",
X"EB",
X"ED",
X"F2",
X"E4",
X"E5",
X"EB",
X"F0",
X"E3",
X"E0",
X"FA",
X"01",
X"04",
X"08",
X"0B",
X"0F",
X"01",
X"FE",
X"05",
X"1A",
X"22",
X"20",
X"34",
X"3E",
X"3E",
X"40",
X"40",
X"43",
X"33",
X"1F",
X"09",
X"03",
X"01",
X"FC",
X"03",
X"0D",
X"06",
X"04",
X"00",
X"FD",
X"FA",
X"E8",
X"E7",
X"E9",
X"E9",
X"EA",
X"EB",
X"EC",
X"ED",
X"EE",
X"EF",
X"EF",
X"F0",
X"F1",
X"F1",
X"F2",
X"F3",
X"F3",
X"F4",
X"F4",
X"F5",
X"F5",
X"F6",
X"F6",
X"F7",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"08",
X"1D",
X"16",
X"14",
X"17",
X"0E",
X"09",
X"0C",
X"19",
X"19",
X"0E",
X"11",
X"15",
X"04",
X"0E",
X"10",
X"06",
X"0C",
X"0F",
X"05",
X"0A",
X"1D",
X"02",
X"F4",
X"13",
X"F8",
X"F5",
X"F7",
X"FE",
X"FB",
X"EF",
X"E8",
X"EB",
X"DF",
X"C9",
X"CC",
X"DE",
X"EE",
X"F7",
X"01",
X"1B",
X"1F",
X"0C",
X"19",
X"1C",
X"2B",
X"20",
X"23",
X"04",
X"01",
X"03",
X"F4",
X"E5",
X"E2",
X"E0",
X"DF",
X"DB",
X"D4",
X"F8",
X"F4",
X"FF",
X"0A",
X"09",
X"1A",
X"2A",
X"34",
X"31",
X"28",
X"1F",
X"1F",
X"FC",
X"F0",
X"E6",
X"DC",
X"E5",
X"DA",
X"C8",
X"D5",
X"E7",
X"F2",
X"F5",
X"08",
X"17",
X"26",
X"2E",
X"23",
X"39",
X"2C",
X"10",
X"16",
X"0E",
X"EB",
X"F2",
X"E7",
X"D9",
X"D3",
X"DC",
X"E9",
X"D5",
X"E5",
X"F4",
X"F7",
X"06",
X"1D",
X"1E",
X"21",
X"33",
X"33",
X"29",
X"1C",
X"05",
X"0B",
X"F5",
X"E0",
X"F2",
X"D1",
X"BE",
X"D1",
X"CE",
X"EE",
X"ED",
X"02",
X"07",
X"11",
X"1E",
X"25",
X"2D",
X"34",
X"2A",
X"28",
X"2B",
X"4E",
X"4C",
X"37",
X"2D",
X"2E",
X"01",
X"B6",
X"BC",
X"DD",
X"D9",
X"E6",
X"1E",
X"1E",
X"3C",
X"6A",
X"62",
X"47",
X"42",
X"2B",
X"1F",
X"1A",
X"27",
X"FE",
X"00",
X"EB",
X"EA",
X"B6",
X"B6",
X"B7",
X"D5",
X"F9",
X"2D",
X"3F",
X"47",
X"56",
X"5F",
X"51",
X"37",
X"F5",
X"FD",
X"DA",
X"F8",
X"01",
X"FC",
X"EE",
X"E6",
X"F3",
X"D3",
X"E0",
X"EE",
X"F7",
X"10",
X"3D",
X"44",
X"25",
X"28",
X"26",
X"F7",
X"05",
X"EA",
X"F1",
X"E8",
X"1C",
X"2D",
X"21",
X"0B",
X"09",
X"E1",
X"C3",
X"DA",
X"D9",
X"B8",
X"F9",
X"03",
X"23",
X"12",
X"2C",
X"08",
X"1A",
X"33",
X"13",
X"07",
X"24",
X"22",
X"17",
X"0A",
X"01",
X"B6",
X"A1",
X"AE",
X"C4",
X"C6",
X"E5",
X"12",
X"1A",
X"3E",
X"53",
X"4C",
X"22",
X"29",
X"25",
X"18",
X"0E",
X"FB",
X"F2",
X"E7",
X"EE",
X"CF",
X"9D",
X"A7",
X"B1",
X"F1",
X"00",
X"3A",
X"34",
X"3C",
X"45",
X"53",
X"33",
X"09",
X"E9",
X"ED",
X"D7",
X"F6",
X"F8",
X"F6",
X"ED",
X"00",
X"E3",
X"D2",
X"DD",
X"E4",
X"FD",
X"10",
X"10",
X"20",
X"FA",
X"1D",
X"06",
X"00",
X"F6",
X"F5",
X"E1",
X"F4",
X"2D",
X"08",
X"11",
X"00",
X"FA",
X"C5",
X"D9",
X"CF",
X"C9",
X"D5",
X"00",
X"0A",
X"1C",
X"26",
X"25",
X"17",
X"1F",
X"12",
X"14",
X"01",
X"21",
X"16",
X"1C",
X"0F",
X"CF",
X"A1",
X"93",
X"B2",
X"BE",
X"BE",
X"EE",
X"0A",
X"45",
X"3F",
X"4E",
X"45",
X"38",
X"17",
X"1C",
X"0A",
X"E6",
X"00",
X"E6",
X"E5",
X"DF",
X"D2",
X"A6",
X"B4",
X"DC",
X"FD",
X"04",
X"33",
X"2D",
X"3C",
X"46",
X"53",
X"16",
X"14",
X"F2",
X"E8",
X"E6",
X"F6",
X"FB",
X"E9",
X"07",
X"01",
X"D2",
X"D4",
X"D5",
X"FB",
X"F7",
X"13",
X"1B",
X"01",
X"1D",
X"2E",
X"14",
X"00",
X"00",
X"F3",
X"FB",
X"20",
X"2A",
X"1A",
X"08",
X"FE",
X"EE",
X"D3",
X"D8",
X"9F",
X"CF",
X"D6",
X"02",
X"00",
X"15",
X"1A",
X"27",
X"35",
X"25",
X"26",
X"12",
X"FD",
X"2B",
X"19",
X"15",
X"DC",
X"D6",
X"C1",
X"AA",
X"AB",
X"CE",
X"C2",
X"F8",
X"2A",
X"3D",
X"36",
X"50",
X"3D",
X"2C",
X"26",
X"1F",
X"FB",
X"F4",
X"FB",
X"D9",
X"E2",
X"D4",
X"CC",
X"99",
X"CB",
X"E1",
X"F3",
X"00",
X"26",
X"3B",
X"3F",
X"2C",
X"2D",
X"F7",
X"05",
X"FF",
X"F2",
X"DE",
X"EF",
X"EA",
X"F8",
X"00",
X"F9",
X"D1",
X"EA",
X"E0",
X"DE",
X"F4",
X"06",
X"FF",
X"07",
X"24",
X"1C",
X"0F",
X"09",
X"00",
X"00",
X"0D",
X"22",
X"23",
X"15",
X"FF",
X"04",
X"DE",
X"CF",
X"AB",
X"C2",
X"CF",
X"E4",
X"0E",
X"10",
X"17",
X"2C",
X"3F",
X"28",
X"28",
X"20",
X"1E",
X"18",
X"1A",
X"08",
X"EF",
X"D1",
X"DE",
X"B4",
X"A2",
X"B6",
X"C9",
X"CF",
X"11",
X"2D",
X"36",
X"37",
X"55",
X"29",
X"29",
X"23",
X"13",
X"E5",
X"FD",
X"00",
X"EA",
X"DB",
X"E5",
X"BE",
X"B7",
X"DD",
X"ED",
X"FF",
X"0F",
X"26",
X"25",
X"3E",
X"3A",
X"0F",
X"14",
X"00",
X"F8",
X"00",
X"E2",
X"FF",
X"FE",
X"00",
X"05",
X"EF",
X"CF",
X"DD",
X"D8",
X"EE",
X"00",
X"FE",
X"00",
X"07",
X"1A",
X"30",
X"16",
X"14",
X"FA",
X"21",
X"13",
X"19",
X"13",
X"0F",
X"FE",
X"00",
X"DD",
X"B8",
X"B4",
X"D1",
X"CF",
X"E9",
X"09",
X"0C",
X"0D",
X"33",
X"3A",
X"2A",
X"24",
X"16",
X"15",
X"0F",
X"0D",
X"F9",
X"DC",
X"D9",
X"CB",
X"C4",
X"BB",
X"AA",
X"D7",
X"D7",
X"20",
X"13",
X"39",
X"2A",
X"41",
X"27",
X"23",
X"12",
X"F5",
X"E5",
X"F9",
X"FB",
X"ED",
X"EB",
X"DE",
X"C8",
X"DC",
X"DB",
X"ED",
X"FA",
X"0E",
X"22",
X"30",
X"26",
X"1C",
X"17",
X"12",
X"08",
X"0C",
X"02",
X"ED",
X"ED",
X"FE",
X"FB",
X"F7",
X"E9",
X"BF",
X"CF",
X"E9",
X"EF",
X"DE",
X"05",
X"06",
X"28",
X"26",
X"1C",
X"1A",
X"04",
X"08",
X"16",
X"04",
X"1D",
X"00",
X"0F",
X"00",
X"FA",
X"BA",
X"BA",
X"CC",
X"D4",
X"CE",
X"F7",
X"11",
X"18",
X"2B",
X"35",
X"3B",
X"2B",
X"1A",
X"1B",
X"0B",
X"26",
X"03",
X"EA",
X"E9",
X"DA",
X"D4",
X"B9",
X"BF",
X"BB",
X"E6",
X"0D",
X"21",
X"23",
X"26",
X"39",
X"47",
X"37",
X"27",
X"00",
X"00",
X"E2",
X"02",
X"FB",
X"EC",
X"E3",
X"E0",
X"D6",
X"DB",
X"E7",
X"EB",
X"E9",
X"19",
X"24",
X"24",
X"1E",
X"1E",
X"0F",
X"0E",
X"0B",
X"F8",
X"D7",
X"E2",
X"FF",
X"FC",
X"EE",
X"E8",
X"CF",
X"BA",
X"C8",
X"D6",
X"CD",
X"D6",
X"FE",
X"00",
X"0D",
X"13",
X"1A",
X"02",
X"14",
X"15",
X"07",
X"02",
X"12",
X"04",
X"FF",
X"F5",
X"DD",
X"A3",
X"AF",
X"BA",
X"CB",
X"D5",
X"FD",
X"03",
X"18",
X"38",
X"3E",
X"2F",
X"26",
X"1D",
X"14",
X"05",
X"0A",
X"F5",
X"EB",
X"DF",
X"DA",
X"BD",
X"AE",
X"BC",
X"CD",
X"F1",
X"09",
X"23",
X"28",
X"32",
X"3B",
X"39",
X"27",
X"0D",
X"FA",
X"F4",
X"EF",
X"00",
X"F0",
X"EC",
X"E0",
X"EA",
X"D0",
X"D6",
X"E0",
X"ED",
X"F9",
X"1C",
X"25",
X"1A",
X"17",
X"25",
X"10",
X"0F",
X"00",
X"FD",
X"EC",
X"0D",
X"18",
X"09",
X"00",
X"F9",
X"DA",
X"CB",
X"DC",
X"D8",
X"D0",
X"F2",
X"07",
X"0F",
X"18",
X"25",
X"1D",
X"1A",
X"2A",
X"19",
X"0F",
X"0D",
X"1B",
X"08",
X"04",
X"F3",
X"CC",
X"AD",
X"B9",
X"C4",
X"D1",
X"E2",
X"05",
X"11",
X"36",
X"3C",
X"43",
X"2E",
X"2C",
X"1B",
X"13",
X"04",
X"FD",
X"F3",
X"ED",
X"E1",
X"DC",
X"BA",
X"B4",
X"C2",
X"E7",
X"F6",
X"09",
X"1D",
X"23",
X"2C",
X"36",
X"32",
X"15",
X"06",
X"00",
X"F2",
X"F4",
X"FA",
X"EF",
X"E4",
X"EC",
X"E6",
X"C8",
X"D6",
X"DF",
X"ED",
X"FA",
X"1B",
X"13",
X"12",
X"1D",
X"23",
X"15",
X"12",
X"05",
X"FC",
X"FC",
X"18",
X"09",
X"01",
X"F6",
X"F1",
X"CF",
X"D0",
X"D4",
X"CF",
X"DB",
X"FA",
X"09",
X"11",
X"1A",
X"24",
X"22",
X"2E",
X"24",
X"19",
X"0B",
X"0E",
X"10",
X"03",
X"F9",
X"DC",
X"C8",
X"B3",
X"C0",
X"CD",
X"D8",
X"EB",
X"08",
X"22",
X"31",
X"37",
X"3D",
X"2D",
X"2B",
X"1A",
X"12",
X"F6",
X"FC",
X"F3",
X"EA",
X"DF",
X"D8",
X"BB",
X"BB",
X"D8",
X"EF",
X"F5",
X"14",
X"20",
X"2B",
X"2F",
X"3E",
X"24",
X"12",
X"0B",
X"00",
X"F6",
X"FA",
X"FD",
X"EE",
X"F1",
X"F8",
X"DF",
X"CD",
X"D8",
X"E6",
X"EE",
X"03",
X"15",
X"0A",
X"18",
X"1F",
X"24",
X"16",
X"14",
X"04",
X"02",
X"0C",
X"16",
X"09",
X"00",
X"F6",
X"EC",
X"CE",
X"CF",
X"C6",
X"D5",
X"DF",
X"00",
X"0A",
X"15",
X"1C",
X"29",
X"32",
X"2F",
X"21",
X"18",
X"09",
X"10",
X"0D",
X"02",
X"E5",
X"DA",
X"C4",
X"B5",
X"C4",
X"D0",
X"DB",
X"F0",
X"1B",
X"28",
X"30",
X"3B",
X"39",
X"2D",
X"26",
X"1B",
X"00",
X"F1",
X"FF",
X"F0",
X"EB",
X"DE",
X"D6",
X"B5",
X"CB",
X"E3",
X"EE",
X"FA",
X"17",
X"22",
X"2B",
X"35",
X"33",
X"16",
X"15",
X"06",
X"00",
X"F2",
X"FF",
X"F7",
X"F6",
X"FC",
X"F4",
X"DA",
X"CE",
X"DC",
X"E7",
X"F1",
X"03",
X"07",
X"0E",
X"17",
X"22",
X"21",
X"16",
X"10",
X"07",
X"10",
X"0D",
X"15",
X"06",
X"00",
X"F5",
X"E8",
X"CA",
X"C0",
X"C7",
X"D7",
X"E2",
X"04",
X"0B",
X"17",
X"1D",
X"3A",
X"32",
X"2D",
X"20",
X"15",
X"08",
X"12",
X"0C",
X"F3",
X"DE",
X"DD",
X"BD",
X"B9",
X"C4",
X"D4",
X"DA",
X"03",
X"24",
X"27",
X"31",
X"3C",
X"38",
X"2B",
X"26",
X"0F",
X"F4",
X"F7",
X"FC",
X"F1",
X"E6",
X"E0",
X"CE",
X"BE",
X"DA",
X"E3",
X"F0",
X"FD",
X"1C",
X"22",
X"2D",
X"2E",
X"23",
X"18",
X"13",
X"07",
X"FF",
X"F4",
X"FF",
X"FA",
X"03",
X"F9",
X"F1",
X"D4",
X"CF",
X"DD",
X"E8",
X"ED",
X"D9",
X"D9",
X"DB",
X"DC",
X"DE",
X"E0",
X"E1",
X"E2",
X"E3",
X"E5",
X"E6",
X"E7",
X"E8",
X"E9",
X"EA",
X"EB",
X"EC",
X"ED",
X"ED",
X"EE",
X"EF",
X"F0",
X"F0",
X"F1",
X"F2",
X"F3",
X"F3",
X"F4",
X"F4",
X"F5",
X"F5",
X"F6",
X"F6",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"07",
X"11",
X"14",
X"14",
X"22",
X"1B",
X"09",
X"0D",
X"00",
X"03",
X"08",
X"0C",
X"07",
X"08",
X"17",
X"1A",
X"11",
X"F1",
X"0C",
X"00",
X"04",
X"FB",
X"07",
X"06",
X"06",
X"04",
X"00",
X"15",
X"09",
X"02",
X"01",
X"02",
X"0D",
X"07",
X"06",
X"0F",
X"01",
X"08",
X"0B",
X"07",
X"00",
X"04",
X"03",
X"0A",
X"00",
X"FF",
X"0D",
X"03",
X"03",
X"0F",
X"0F",
X"F6",
X"05",
X"00",
X"F3",
X"08",
X"FA",
X"03",
X"FB",
X"09",
X"02",
X"10",
X"F8",
X"FE",
X"06",
X"02",
X"F2",
X"FD",
X"FF",
X"06",
X"00",
X"01",
X"06",
X"10",
X"FD",
X"FD",
X"03",
X"F9",
X"02",
X"14",
X"F1",
X"F9",
X"FF",
X"F7",
X"06",
X"ED",
X"FF",
X"F5",
X"05",
X"F9",
X"FE",
X"06",
X"0C",
X"F5",
X"04",
X"0A",
X"FE",
X"05",
X"03",
X"06",
X"08",
X"0B",
X"F3",
X"FB",
X"00",
X"00",
X"00",
X"FC",
X"05",
X"FC",
X"FD",
X"04",
X"0E",
X"0F",
X"F9",
X"F6",
X"FC",
X"F5",
X"0C",
X"FE",
X"FE",
X"F4",
X"FE",
X"FF",
X"10",
X"01",
X"FA",
X"0D",
X"00",
X"E8",
X"03",
X"F0",
X"FC",
X"F4",
X"06",
X"02",
X"FF",
X"FF",
X"01",
X"00",
X"FE",
X"0B",
X"00",
X"09",
X"0F",
X"FB",
X"F9",
X"05",
X"F7",
X"F6",
X"01",
X"03",
X"F6",
X"02",
X"00",
X"09",
X"0C",
X"00",
X"FC",
X"03",
X"F3",
X"09",
X"06",
X"FC",
X"F9",
X"F9",
X"07",
X"0E",
X"E6",
X"03",
X"F3",
X"FF",
X"00",
X"FF",
X"06",
X"F8",
X"F6",
X"02",
X"04",
X"FB",
X"FF",
X"02",
X"04",
X"0A",
X"01",
X"F8",
X"05",
X"00",
X"01",
X"FE",
X"00",
X"FD",
X"FF",
X"08",
X"07",
X"01",
X"09",
X"FB",
X"00",
X"07",
X"05",
X"01",
X"F6",
X"FA",
X"FC",
X"F7",
X"FD",
X"FE",
X"05",
X"04",
X"0A",
X"F9",
X"FE",
X"FF",
X"03",
X"05",
X"F8",
X"05",
X"F7",
X"FE",
X"08",
X"00",
X"00",
X"05",
X"04",
X"08",
X"02",
X"F7",
X"ED",
X"FA",
X"FE",
X"FE",
X"FC",
X"00",
X"06",
X"01",
X"FF",
X"FF",
X"03",
X"00",
X"09",
X"FD",
X"F6",
X"04",
X"FE",
X"FD",
X"FB",
X"05",
X"00",
X"05",
X"0B",
X"EF",
X"03",
X"06",
X"F0",
X"FA",
X"F9",
X"FF",
X"FF",
X"04",
X"06",
X"01",
X"07",
X"F9",
X"F4",
X"FB",
X"00",
X"06",
X"FF",
X"03",
X"05",
X"00",
X"FA",
X"0D",
X"0B",
X"FB",
X"FB",
X"04",
X"F6",
X"FF",
X"09",
X"FA",
X"FB",
X"07",
X"04",
X"03",
X"FF",
X"00",
X"FE",
X"00",
X"FF",
X"01",
X"09",
X"02",
X"FB",
X"05",
X"04",
X"00",
X"05",
X"09",
X"EC",
X"F4",
X"FF",
X"F6",
X"00",
X"F5",
X"0D",
X"FB",
X"FF",
X"F4",
X"FF",
X"00",
X"09",
X"08",
X"FB",
X"07",
X"09",
X"E9",
X"07",
X"FA",
X"FD",
X"F9",
X"06",
X"0A",
X"01",
X"FA",
X"FD",
X"F7",
X"09",
X"FB",
X"FA",
X"FE",
X"00",
X"10",
X"05",
X"00",
X"F6",
X"F2",
X"F5",
X"FD",
X"FD",
X"FC",
X"00",
X"0D",
X"10",
X"F9",
X"F4",
X"02",
X"EE",
X"02",
X"00",
X"00",
X"F6",
X"00",
X"00",
X"08",
X"FC",
X"05",
X"0E",
X"FE",
X"FD",
X"06",
X"F9",
X"00",
X"0A",
X"05",
X"FB",
X"03",
X"00",
X"00",
X"FE",
X"02",
X"05",
X"F9",
X"FD",
X"08",
X"07",
X"FE",
X"08",
X"00",
X"EE",
X"07",
X"FD",
X"05",
X"FA",
X"F4",
X"07",
X"FF",
X"05",
X"F5",
X"00",
X"0D",
X"F9",
X"FD",
X"F8",
X"FB",
X"0B",
X"FC",
X"06",
X"FB",
X"00",
X"09",
X"0B",
X"00",
X"FB",
X"00",
X"FD",
X"0F",
X"03",
X"F4",
X"FB",
X"F3",
X"09",
X"00",
X"00",
X"FB",
X"F5",
X"04",
X"00",
X"03",
X"FF",
X"00",
X"08",
X"06",
X"02",
X"FF",
X"F9",
X"F7",
X"07",
X"0B",
X"E8",
X"FE",
X"F6",
X"06",
X"03",
X"E9",
X"00",
X"F6",
X"F8",
X"F9",
X"01",
X"03",
X"00",
X"FB",
X"05",
X"0D",
X"FA",
X"FC",
X"02",
X"00",
X"0C",
X"00",
X"F4",
X"FE",
X"00",
X"03",
X"FA",
X"00",
X"05",
X"00",
X"00",
X"07",
X"0A",
X"0D",
X"F9",
X"00",
X"F6",
X"00",
X"06",
X"F8",
X"00",
X"F6",
X"03",
X"0D",
X"F1",
X"02",
X"00",
X"FF",
X"05",
X"FF",
X"01",
X"FD",
X"FB",
X"01",
X"0B",
X"06",
X"07",
X"FA",
X"00",
X"FC",
X"0A",
X"0F",
X"F8",
X"F2",
X"FF",
X"F1",
X"FF",
X"00",
X"00",
X"F4",
X"03",
X"03",
X"04",
X"FB",
X"02",
X"0D",
X"0C",
X"F3",
X"00",
X"F2",
X"F5",
X"FA",
X"FC",
X"00",
X"FB",
X"0C",
X"03",
X"02",
X"E9",
X"00",
X"FB",
X"FE",
X"FD",
X"FF",
X"09",
X"05",
X"02",
X"F2",
X"01",
X"02",
X"0E",
X"04",
X"EA",
X"0B",
X"F6",
X"00",
X"FC",
X"04",
X"00",
X"00",
X"08",
X"F4",
X"00",
X"00",
X"03",
X"05",
X"F4",
X"00",
X"01",
X"01",
X"05",
X"0C",
X"02",
X"01",
X"EF",
X"FD",
X"FB",
X"FF",
X"F9",
X"04",
X"07",
X"0C",
X"FF",
X"F3",
X"08",
X"FD",
X"02",
X"EE",
X"F7",
X"FD",
X"00",
X"FC",
X"00",
X"0D",
X"0E",
X"00",
X"F9",
X"F8",
X"FB",
X"05",
X"0F",
X"FE",
X"FC",
X"01",
X"FE",
X"05",
X"0A",
X"FB",
X"FF",
X"0B",
X"FF",
X"FA",
X"0E",
X"FC",
X"F9",
X"0F",
X"FD",
X"FA",
X"00",
X"FD",
X"01",
X"01",
X"04",
X"FD",
X"FA",
X"0A",
X"0A",
X"FC",
X"FE",
X"00",
X"F7",
X"05",
X"0E",
X"F5",
X"FC",
X"00",
X"F9",
X"00",
X"08",
X"05",
X"F7",
X"09",
X"FF",
X"F8",
X"02",
X"08",
X"F9",
X"00",
X"02",
X"F6",
X"FD",
X"F8",
X"FF",
X"01",
X"FF",
X"05",
X"00",
X"06",
X"0D",
X"FC",
X"FC",
X"00",
X"FA",
X"FF",
X"0C",
X"0C",
X"F6",
X"F8",
X"F7",
X"F9",
X"06",
X"04",
X"03",
X"F0",
X"00",
X"FD",
X"00",
X"03",
X"00",
X"0B",
X"FC",
X"FA",
X"08",
X"00",
X"EE",
X"E8",
X"EB",
X"EB",
X"EC",
X"EC",
X"EE",
X"EF",
X"F0",
X"F0",
X"F1",
X"F1",
X"F3",
X"F4",
X"F4",
X"F4",
X"F5",
X"F4",
X"F5",
X"F6",
X"F7",
X"F7",
X"F6",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FE",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"04",
X"09",
X"0D",
X"12",
X"16",
X"1A",
X"1E",
X"22",
X"26",
X"29",
X"2D",
X"30",
X"33",
X"35",
X"34",
X"2F",
X"27",
X"20",
X"19",
X"13",
X"0D",
X"07",
X"02",
X"FF",
X"FA",
X"F5",
X"F0",
X"EC",
X"E7",
X"E3",
X"E0",
X"DC",
X"D9",
X"D5",
X"D4",
X"D7",
X"DE",
X"E4",
X"EB",
X"F1",
X"F7",
X"FC",
X"00",
X"04",
X"09",
X"0E",
X"12",
X"17",
X"1B",
X"1F",
X"23",
X"26",
X"2A",
X"2D",
X"30",
X"2E",
X"29",
X"21",
X"1B",
X"14",
X"0E",
X"08",
X"03",
X"00",
X"FB",
X"F6",
X"F1",
X"EC",
X"E8",
X"E4",
X"E0",
X"DD",
X"D9",
X"D5",
X"D2",
X"D1",
X"D5",
X"DC",
X"E3",
X"E9",
X"EF",
X"F4",
X"FB",
X"00",
X"02",
X"07",
X"0C",
X"11",
X"15",
X"1A",
X"1F",
X"21",
X"25",
X"29",
X"2C",
X"30",
X"2E",
X"28",
X"20",
X"19",
X"13",
X"30",
X"3A",
X"0C",
X"F7",
X"F7",
X"F0",
X"EE",
X"E7",
X"E5",
X"DE",
X"DF",
X"D5",
X"EB",
X"02",
X"F8",
X"FA",
X"F9",
X"00",
X"02",
X"0A",
X"0B",
X"16",
X"0A",
X"ED",
X"F6",
X"FA",
X"00",
X"02",
X"08",
X"0C",
X"12",
X"14",
X"1D",
X"48",
X"4E",
X"4E",
X"4C",
X"44",
X"3D",
X"33",
X"2D",
X"25",
X"20",
X"F8",
X"E4",
X"E5",
X"DD",
X"DD",
X"D6",
X"D5",
X"CE",
X"D0",
X"C7",
X"E1",
X"F7",
X"EC",
X"EE",
X"EE",
X"F7",
X"F9",
X"00",
X"01",
X"0C",
X"00",
X"E3",
X"EE",
X"F1",
X"F9",
X"FD",
X"02",
X"05",
X"0B",
X"0D",
X"1A",
X"44",
X"48",
X"49",
X"45",
X"3D",
X"35",
X"2E",
X"28",
X"21",
X"1B",
X"F0",
X"E1",
X"E1",
X"DA",
X"D9",
X"D3",
X"D3",
X"CC",
X"CD",
X"C4",
X"E2",
X"F4",
X"EA",
X"ED",
X"EE",
X"F7",
X"F9",
X"00",
X"01",
X"0C",
X"FC",
X"E2",
X"EE",
X"F0",
X"F8",
X"FB",
X"01",
X"04",
X"0C",
X"0C",
X"1C",
X"46",
X"47",
X"49",
X"44",
X"3D",
X"34",
X"2D",
X"27",
X"20",
X"18",
X"EB",
X"E0",
X"DF",
X"DA",
X"D8",
X"D3",
X"D2",
X"CD",
X"CC",
X"C5",
X"E2",
X"EE",
X"E4",
X"E7",
X"E9",
X"F2",
X"F5",
X"FD",
X"FE",
X"08",
X"F8",
X"E4",
X"F0",
X"F2",
X"FA",
X"FD",
X"02",
X"06",
X"0E",
X"0E",
X"20",
X"43",
X"42",
X"45",
X"40",
X"39",
X"30",
X"2A",
X"22",
X"1C",
X"11",
X"EA",
X"E4",
X"E1",
X"DC",
X"DA",
X"D5",
X"D3",
X"CE",
X"CD",
X"C9",
X"E7",
X"EE",
X"E6",
X"E9",
X"EB",
X"F4",
X"F7",
X"FF",
X"00",
X"09",
X"F5",
X"E6",
X"F2",
X"F4",
X"FC",
X"FE",
X"05",
X"07",
X"0F",
X"0F",
X"24",
X"45",
X"42",
X"45",
X"3E",
X"39",
X"2F",
X"29",
X"21",
X"1D",
X"0F",
X"E9",
X"E5",
X"E1",
X"DE",
X"DA",
X"D6",
X"D3",
X"CF",
X"CD",
X"CA",
X"E9",
X"ED",
X"E6",
X"E9",
X"ED",
X"F4",
X"F8",
X"00",
X"00",
X"0A",
X"F3",
X"E7",
X"F2",
X"F4",
X"FD",
X"FF",
X"05",
X"07",
X"10",
X"0E",
X"28",
X"46",
X"43",
X"46",
X"3E",
X"39",
X"2F",
X"29",
X"20",
X"1E",
X"0C",
X"E7",
X"E5",
X"DF",
X"DD",
X"D9",
X"D6",
X"D2",
X"D0",
X"CC",
X"CC",
X"EC",
X"EC",
X"E7",
X"E9",
X"ED",
X"F5",
X"F9",
X"00",
X"FF",
X"03",
X"EE",
X"E9",
X"F3",
X"F5",
X"FE",
X"00",
X"06",
X"09",
X"11",
X"10",
X"2A",
X"41",
X"3F",
X"41",
X"3A",
X"33",
X"2A",
X"25",
X"1B",
X"19",
X"06",
X"E8",
X"E7",
X"E1",
X"DF",
X"DA",
X"D7",
X"D3",
X"D1",
X"CC",
X"CE",
X"E9",
X"E6",
X"E3",
X"E5",
X"EA",
X"F1",
X"F6",
X"FC",
X"00",
X"05",
X"EF",
X"ED",
X"F5",
X"F9",
X"00",
X"02",
X"09",
X"0C",
X"13",
X"13",
X"2F",
X"42",
X"40",
X"42",
X"3A",
X"34",
X"2A",
X"25",
X"1C",
X"1A",
X"03",
X"E8",
X"E8",
X"E2",
X"E0",
X"DA",
X"D8",
X"D3",
X"D2",
X"CC",
X"D1",
X"EA",
X"E5",
X"E3",
X"E5",
X"EC",
X"F2",
X"F7",
X"FD",
X"00",
X"04",
X"EE",
X"EE",
X"F6",
X"FA",
X"00",
X"03",
X"09",
X"0C",
X"13",
X"14",
X"31",
X"42",
X"40",
X"42",
X"39",
X"33",
X"2A",
X"25",
X"1B",
X"1A",
X"01",
X"E8",
X"E9",
X"E2",
X"E0",
X"DA",
X"D8",
X"D3",
X"D2",
X"CC",
X"D4",
X"EB",
X"E5",
X"E4",
X"E5",
X"EC",
X"F2",
X"F8",
X"FD",
X"01",
X"03",
X"EC",
X"EF",
X"F6",
X"FB",
X"00",
X"04",
X"09",
X"0D",
X"13",
X"15",
X"30",
X"3C",
X"3C",
X"3C",
X"34",
X"2D",
X"25",
X"20",
X"17",
X"15",
X"FE",
X"EA",
X"EA",
X"E3",
X"E1",
X"DC",
X"DA",
X"D5",
X"D4",
X"CD",
X"D6",
X"E8",
X"E0",
X"E0",
X"E2",
X"EA",
X"EF",
X"F5",
X"FA",
X"00",
X"00",
X"EE",
X"F3",
X"F9",
X"FE",
X"02",
X"07",
X"0C",
X"10",
X"15",
X"19",
X"35",
X"3E",
X"3E",
X"3D",
X"35",
X"2E",
X"26",
X"21",
X"18",
X"15",
X"FD",
X"EB",
X"EB",
X"E4",
X"E2",
X"DD",
X"DB",
X"D5",
X"D5",
X"CD",
X"D9",
X"E9",
X"E1",
X"E1",
X"E3",
X"EB",
X"EF",
X"F7",
X"FA",
X"00",
X"00",
X"ED",
X"F4",
X"F9",
X"FF",
X"02",
X"08",
X"0C",
X"11",
X"15",
X"1B",
X"37",
X"3E",
X"3E",
X"3C",
X"35",
X"2E",
X"26",
X"20",
X"18",
X"14",
X"FA",
X"EB",
X"EA",
X"E4",
X"E2",
X"DC",
X"DA",
X"D5",
X"D4",
X"CD",
X"DB",
X"E9",
X"E1",
X"E2",
X"E4",
X"EC",
X"F0",
X"F8",
X"FB",
X"02",
X"FE",
X"ED",
X"F6",
X"FA",
X"00",
X"02",
X"08",
X"0C",
X"11",
X"14",
X"1D",
X"39",
X"3E",
X"3F",
X"3C",
X"34",
X"2D",
X"26",
X"20",
X"18",
X"13",
X"F7",
X"EB",
X"E9",
X"E3",
X"E1",
X"DC",
X"DA",
X"D5",
X"D3",
X"CD",
X"DD",
X"E8",
X"E0",
X"E2",
X"E5",
X"ED",
X"F1",
X"F9",
X"FC",
X"03",
X"FC",
X"ED",
X"F7",
X"FA",
X"00",
X"03",
X"09",
X"0C",
X"12",
X"14",
X"1F",
X"3B",
X"3D",
X"3F",
X"3B",
X"34",
X"2C",
X"25",
X"1E",
X"18",
X"11",
X"F5",
X"EB",
X"E9",
X"E3",
X"E1",
X"DC",
X"D9",
X"D4",
X"D3",
X"CD",
X"DF",
X"E8",
X"E0",
X"E2",
X"E4",
X"ED",
X"F1",
X"F9",
X"FC",
X"03",
X"FA",
X"EE",
X"F7",
X"FB",
X"00",
X"03",
X"0A",
X"0D",
X"14",
X"15",
X"22",
X"3C",
X"3D",
X"3F",
X"3A",
X"33",
X"2B",
X"25",
X"1D",
X"18",
X"0F",
X"F3",
X"EB",
X"E8",
X"E3",
X"E0",
X"DC",
X"D9",
X"D5",
X"D3",
X"CD",
X"E1",
X"E7",
X"E0",
X"E2",
X"E5",
X"EE",
X"F2",
X"FA",
X"FC",
X"03",
X"F9",
X"EE",
X"F8",
X"FB",
X"01",
X"04",
X"0A",
X"0D",
X"14",
X"14",
X"24",
X"3D",
X"3D",
X"3F",
X"39",
X"32",
X"2A",
X"24",
X"1D",
X"18",
X"0D",
X"F1",
X"EC",
X"E8",
X"E4",
X"E0",
X"DC",
X"D8",
X"D4",
X"D2",
X"CE",
X"DE",
X"E0",
X"DB",
X"DD",
X"E1",
X"E9",
X"EE",
X"F5",
X"F9",
X"00",
X"F6",
X"F1",
X"FA",
X"FE",
X"02",
X"06",
X"0C",
X"0F",
X"16",
X"16",
X"26",
X"39",
X"39",
X"3B",
X"35",
X"2F",
X"26",
X"21",
X"19",
X"14",
X"09",
X"F2",
X"EF",
X"EA",
X"E6",
X"E2",
X"DE",
X"DA",
X"D6",
X"D3",
X"D1",
X"E2",
X"E1",
X"DC",
X"DE",
X"E3",
X"EB",
X"F0",
X"F7",
X"FB",
X"00",
X"F6",
X"F3",
X"FC",
X"FF",
X"04",
X"07",
X"0D",
X"11",
X"17",
X"18",
X"29",
X"3A",
X"3A",
X"3B",
X"35",
X"2F",
X"26",
X"21",
X"19",
X"15",
X"07",
X"F2",
X"EF",
X"E9",
X"E6",
X"E1",
X"DE",
X"DA",
X"D7",
X"D3",
X"D2",
X"E3",
X"E0",
X"DD",
X"DF",
X"E4",
X"EB",
X"F1",
X"F8",
X"FC",
X"01",
X"F5",
X"F4",
X"FC",
X"00",
X"04",
X"08",
X"0E",
X"11",
X"17",
X"18",
X"2B",
X"3B",
X"3A",
X"3C",
X"35",
X"2E",
X"26",
X"21",
X"18",
X"15",
X"05",
X"F1",
X"EE",
X"E8",
X"E5",
X"E1",
X"DD",
X"D9",
X"D7",
X"D2",
X"D4",
X"E4",
X"DF",
X"DD",
X"E0",
X"E6",
X"ED",
X"F2",
X"F8",
X"FD",
X"00",
X"F4",
X"F5",
X"FC",
X"00",
X"04",
X"08",
X"0E",
X"11",
X"17",
X"19",
X"2D",
X"3A",
X"3A",
X"3B",
X"34",
X"2E",
X"25",
X"20",
X"18",
X"15",
X"03",
X"F0",
X"EF",
X"E8",
X"E6",
X"E0",
X"DE",
X"D9",
X"D7",
X"D1",
X"D5",
X"E4",
X"DE",
X"DD",
X"DF",
X"E6",
X"EC",
X"F3",
X"F8",
X"FE",
X"00",
X"F3",
X"F6",
X"FD",
X"00",
X"05",
X"09",
X"0F",
X"12",
X"18",
X"1A",
X"30",
X"3B",
X"3A",
X"3B",
X"33",
X"2D",
X"25",
X"1F",
X"17",
X"14",
X"00",
X"F0",
X"EE",
X"E8",
X"E5",
X"E0",
X"DD",
X"D9",
X"D7",
X"D1",
X"D6",
X"E4",
X"DE",
X"DE",
X"E0",
X"E7",
X"ED",
X"F3",
X"F8",
X"FF",
X"00",
X"F3",
X"F8",
X"FE",
X"00",
X"05",
X"0A",
X"0E",
X"13",
X"17",
X"1B",
X"31",
X"3A",
X"3A",
X"3A",
X"32",
X"2C",
X"24",
X"1E",
X"16",
X"13",
X"00",
X"EF",
X"EE",
X"E7",
X"E5",
X"E0",
X"DD",
X"D8",
X"D7",
X"D0",
X"D8",
X"E5",
X"DD",
X"DE",
X"E0",
X"E8",
X"ED",
X"F4",
X"F8",
X"00",
X"FF",
X"F2",
X"F7",
X"FD",
X"00",
X"05",
X"0A",
X"0F",
X"12",
X"11",
X"11",
X"10",
X"0F",
X"0E",
X"0E",
X"0D",
X"0C",
X"0C",
X"0B",
X"0B",
X"0A",
X"0A",
X"09",
X"09",
X"08",
X"08",
X"08",
X"07",
X"07",
X"07",
X"06",
X"06",
X"05",
X"05",
X"05",
X"05",
X"04",
X"04",
X"04",
X"04",
X"03",
X"03",
X"03",
X"03",
X"03",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"02",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"18",
X"24",
X"0A",
X"10",
X"11",
X"10",
X"1B",
X"03",
X"0D",
X"08",
X"09",
X"14",
X"04",
X"16",
X"08",
X"08",
X"14",
X"0A",
X"0D",
X"0E",
X"05",
X"0A",
X"12",
X"06",
X"FD",
X"06",
X"0C",
X"0C",
X"FF",
X"FF",
X"06",
X"03",
X"0A",
X"0C",
X"15",
X"00",
X"FE",
X"FB",
X"FF",
X"FF",
X"11",
X"06",
X"F9",
X"0A",
X"09",
X"EF",
X"06",
X"02",
X"FC",
X"00",
X"F8",
X"02",
X"03",
X"07",
X"FF",
X"06",
X"06",
X"0A",
X"01",
X"09",
X"00",
X"FF",
X"06",
X"0B",
X"FD",
X"00",
X"F1",
X"FD",
X"FF",
X"FE",
X"FB",
X"03",
X"0C",
X"08",
X"00",
X"FE",
X"00",
X"01",
X"12",
X"04",
X"FD",
X"F8",
X"F9",
X"FC",
X"08",
X"0E",
X"EB",
X"FF",
X"04",
X"F6",
X"F6",
X"F2",
X"F8",
X"00",
X"00",
X"FC",
X"04",
X"08",
X"03",
X"F9",
X"05",
X"07",
X"00",
X"FB",
X"15",
X"00",
X"F0",
X"00",
X"F3",
X"00",
X"FE",
X"07",
X"FB",
X"00",
X"00",
X"FE",
X"0A",
X"FF",
X"07",
X"10",
X"00",
X"F8",
X"07",
X"F5",
X"FE",
X"02",
X"07",
X"EF",
X"00",
X"00",
X"FF",
X"F1",
X"E9",
X"EC",
X"EC",
X"EE",
X"EE",
X"F0",
X"F0",
X"F0",
X"F2",
X"F2",
X"F3",
X"F3",
X"F5",
X"F4",
X"F5",
X"F6",
X"F6",
X"F6",
X"F6",
X"F7",
X"F6",
X"F8",
X"F8",
X"F9",
X"F8",
X"FA",
X"F9",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"13",
X"0C",
X"1A",
X"13",
X"13",
X"18",
X"13",
X"16",
X"1D",
X"07",
X"00",
X"0A",
X"0C",
X"04",
X"00",
X"0F",
X"09",
X"10",
X"07",
X"18",
X"1C",
X"08",
X"EF",
X"04",
X"F1",
X"0F",
X"FE",
X"04",
X"F9",
X"0A",
X"00",
X"04",
X"06",
X"02",
X"0E",
X"02",
X"02",
X"04",
X"0A",
X"FE",
X"00",
X"0B",
X"13",
X"01",
X"06",
X"00",
X"04",
X"0F",
X"12",
X"FF",
X"FE",
X"FA",
X"FE",
X"00",
X"0E",
X"0B",
X"EA",
X"0E",
X"FC",
X"F6",
X"FE",
X"FA",
X"01",
X"FE",
X"03",
X"03",
X"04",
X"FC",
X"0F",
X"00",
X"01",
X"0C",
X"FF",
X"02",
X"12",
X"FF",
X"F1",
X"FF",
X"F5",
X"04",
X"01",
X"00",
X"00",
X"FB",
X"FE",
X"02",
X"06",
X"03",
X"07",
X"07",
X"00",
X"FE",
X"F6",
X"F9",
X"FD",
X"FC",
X"01",
X"FF",
X"0D",
X"05",
X"03",
X"05",
X"F9",
X"FA",
X"0D",
X"FC",
X"FD",
X"03",
X"03",
X"0F",
X"F8",
X"FB",
X"02",
X"F9",
X"00",
X"08",
X"06",
X"FF",
X"07",
X"00",
X"F9",
X"FE",
X"04",
X"06",
X"01",
X"FB",
X"00",
X"00",
X"04",
X"02",
X"04",
X"F2",
X"E7",
X"EB",
X"E8",
X"EC",
X"ED",
X"ED",
X"EE",
X"EF",
X"F1",
X"F0",
X"F1",
X"F2",
X"F2",
X"F3",
X"F3",
X"F4",
X"F5",
X"F5",
X"F6",
X"F6",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"06",
X"18",
X"14",
X"1C",
X"11",
X"08",
X"1A",
X"1B",
X"0B",
X"04",
X"08",
X"0A",
X"13",
X"0C",
X"13",
X"0B",
X"0C",
X"05",
X"0D",
X"10",
X"0B",
X"05",
X"13",
X"00",
X"03",
X"11",
X"0F",
X"F6",
X"00",
X"00",
X"08",
X"F7",
X"00",
X"04",
X"08",
X"09",
X"00",
X"0D",
X"13",
X"03",
X"FB",
X"0B",
X"F4",
X"06",
X"0C",
X"F2",
X"FC",
X"FD",
X"01",
X"0A",
X"FA",
X"00",
X"00",
X"FE",
X"FE",
X"07",
X"04",
X"00",
X"09",
X"0C",
X"09",
X"FA",
X"03",
X"FD",
X"06",
X"0F",
X"00",
X"F5",
X"FF",
X"FA",
X"08",
X"F8",
X"00",
X"FF",
X"F7",
X"00",
X"00",
X"08",
X"09",
X"00",
X"01",
X"01",
X"EF",
X"04",
X"FD",
X"FC",
X"FE",
X"07",
X"16",
X"00",
X"EC",
X"08",
X"E9",
X"FF",
X"F3",
X"00",
X"F0",
X"05",
X"FC",
X"0C",
X"FF",
X"F5",
X"08",
X"FA",
X"00",
X"FD",
X"0C",
X"05",
X"08",
X"01",
X"00",
X"FE",
X"01",
X"06",
X"00",
X"05",
X"07",
X"00",
X"00",
X"07",
X"05",
X"FC",
X"0C",
X"FD",
X"E9",
X"00",
X"F4",
X"03",
X"F4",
X"00",
X"0A",
X"F0",
X"ED",
X"E9",
X"EE",
X"EB",
X"EF",
X"EE",
X"F1",
X"EF",
X"F3",
X"F1",
X"F3",
X"F2",
X"F4",
X"F3",
X"F5",
X"F4",
X"F6",
X"F5",
X"F7",
X"F7",
X"F7",
X"F7",
X"F9",
X"F7",
X"F9",
X"F8",
X"FA",
X"F9",
X"FB",
X"F9",
X"FB",
X"F9",
X"FB",
X"FB",
X"FC",
X"FC",
X"FD",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FD",
X"1D",
X"2E",
X"28",
X"28",
X"25",
X"24",
X"22",
X"FD",
X"F3",
X"F7",
X"F5",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F9",
X"F8",
X"FA",
X"F7",
X"02",
X"28",
X"22",
X"25",
X"FC",
X"F4",
X"F3",
X"05",
X"27",
X"23",
X"2A",
X"00",
X"0A",
X"04",
X"26",
X"31",
X"29",
X"19",
X"EF",
X"EC",
X"E7",
X"E1",
X"E1",
X"D8",
X"EA",
X"03",
X"FC",
X"F9",
X"F2",
X"ED",
X"EC",
X"CB",
X"B0",
X"B4",
X"BA",
X"E9",
X"EA",
X"F7",
X"D6",
X"D0",
X"DA",
X"E0",
X"E8",
X"EC",
X"F4",
X"F7",
X"00",
X"00",
X"1F",
X"3D",
X"38",
X"40",
X"3F",
X"43",
X"42",
X"41",
X"37",
X"30",
X"29",
X"23",
X"1C",
X"16",
X"0F",
X"09",
X"02",
X"00",
X"FC",
X"F7",
X"EC",
X"BF",
X"C1",
X"B7",
X"D9",
X"E5",
X"E2",
X"D3",
X"B3",
X"C3",
X"C6",
X"F7",
X"02",
X"04",
X"0A",
X"0F",
X"14",
X"16",
X"1D",
X"1C",
X"27",
X"07",
X"FC",
X"04",
X"07",
X"0C",
X"12",
X"15",
X"39",
X"3A",
X"33",
X"16",
X"F2",
X"F7",
X"E9",
X"EC",
X"E3",
X"E2",
X"DC",
X"DD",
X"D3",
X"DD",
X"FB",
X"FC",
X"F1",
X"F5",
X"D3",
X"CF",
X"EE",
X"E9",
X"F6",
X"F7",
X"00",
X"00",
X"08",
X"E3",
X"E5",
X"E9",
X"FE",
X"24",
X"26",
X"29",
X"38",
X"61",
X"5C",
X"63",
X"5F",
X"67",
X"61",
X"64",
X"32",
X"EE",
X"EE",
X"E7",
X"E7",
X"DF",
X"DE",
X"DA",
X"FE",
X"00",
X"F9",
X"F5",
X"F2",
X"12",
X"18",
X"FF",
X"D7",
X"D7",
X"D2",
X"D5",
X"DA",
X"E3",
X"E4",
X"09",
X"23",
X"FF",
X"F8",
X"00",
X"04",
X"0A",
X"0B",
X"EB",
X"E9",
X"F1",
X"F7",
X"FE",
X"FF",
X"20",
X"4B",
X"67",
X"60",
X"56",
X"4C",
X"45",
X"3D",
X"37",
X"10",
X"F6",
X"FE",
X"DB",
X"BC",
X"BF",
X"BA",
X"BE",
X"E4",
X"E3",
X"DD",
X"DA",
X"D5",
X"D5",
X"D4",
X"D9",
X"E2",
X"E9",
X"ED",
X"F5",
X"F7",
X"00",
X"00",
X"26",
X"3E",
X"38",
X"41",
X"37",
X"15",
X"1A",
X"19",
X"F7",
X"FC",
X"00",
X"03",
X"FF",
X"FD",
X"F4",
X"02",
X"21",
X"3C",
X"3C",
X"2F",
X"2D",
X"20",
X"1F",
X"F5",
X"E3",
X"E1",
X"DE",
X"D7",
X"D6",
X"AA",
X"A4",
X"D1",
X"D0",
X"D9",
X"DD",
X"E6",
X"E4",
X"F2",
X"DF",
X"CF",
X"D6",
X"F9",
X"10",
X"0C",
X"17",
X"16",
X"3D",
X"49",
X"4B",
X"4B",
X"4F",
X"4E",
X"54",
X"2E",
X"ED",
X"F0",
X"E4",
X"E7",
X"DE",
X"DF",
X"D6",
X"EB",
X"FC",
X"F5",
X"EE",
X"F8",
X"13",
X"06",
X"05",
X"DE",
X"D3",
X"CE",
X"CE",
X"D0",
X"D7",
X"DB",
X"EF",
X"0B",
X"ED",
X"F7",
X"F7",
X"00",
X"00",
X"0C",
X"FA",
X"E8",
X"F2",
X"F6",
X"FE",
X"03",
X"2D",
X"31",
X"56",
X"5D",
X"54",
X"4B",
X"41",
X"39",
X"34",
X"22",
X"FC",
X"FB",
X"D1",
X"C9",
X"C6",
X"C4",
X"BE",
X"D5",
X"E8",
X"DE",
X"DE",
X"D7",
X"D7",
X"D0",
X"F2",
X"E2",
X"DF",
X"EA",
X"EE",
X"F4",
X"FA",
X"FD",
X"0C",
X"32",
X"2E",
X"3B",
X"20",
X"11",
X"19",
X"1E",
X"08",
X"F9",
X"05",
X"04",
X"09",
X"01",
X"00",
X"F8",
X"28",
X"41",
X"35",
X"2E",
X"27",
X"20",
X"1B",
X"08",
X"E4",
X"E6",
X"DC",
X"DF",
X"CC",
X"AC",
X"A9",
X"C4",
X"D6",
X"D3",
X"DD",
X"E2",
X"EA",
X"EE",
X"F4",
X"D2",
X"DE",
X"05",
X"0B",
X"0E",
X"15",
X"15",
X"27",
X"41",
X"3D",
X"43",
X"42",
X"48",
X"44",
X"29",
X"04",
X"F5",
X"F4",
X"EE",
X"EA",
X"E5",
X"E1",
X"E0",
X"FB",
X"F9",
X"F2",
X"05",
X"0D",
X"01",
X"01",
X"ED",
X"D1",
X"D2",
X"CC",
X"CD",
X"D0",
X"D7",
X"DE",
X"E9",
X"EA",
X"F1",
X"F7",
X"FF",
X"01",
X"06",
X"07",
X"F0",
X"F5",
X"FC",
X"FE",
X"12",
X"2E",
X"29",
X"3F",
X"56",
X"4E",
X"4A",
X"40",
X"3B",
X"31",
X"2B",
X"0B",
X"F1",
X"D6",
X"D4",
X"CF",
X"CD",
X"C9",
X"CB",
X"E6",
X"E2",
X"DF",
X"DB",
X"D8",
X"D7",
X"F8",
X"E8",
X"D9",
X"E4",
X"E6",
X"F0",
X"F3",
X"FC",
X"FE",
X"1F",
X"2A",
X"2A",
X"11",
X"11",
X"16",
X"1B",
X"19",
X"00",
X"06",
X"08",
X"10",
X"0B",
X"0B",
X"00",
X"2A",
X"40",
X"32",
X"2E",
X"22",
X"20",
X"15",
X"14",
X"F0",
X"E6",
X"E0",
X"E1",
X"C5",
X"B4",
X"B3",
X"B7",
X"D5",
X"D1",
X"D9",
X"DC",
X"E7",
X"E7",
X"F6",
X"E2",
X"E7",
X"05",
X"04",
X"0D",
X"0D",
X"15",
X"16",
X"39",
X"42",
X"45",
X"44",
X"4B",
X"3F",
X"29",
X"21",
X"FE",
X"FC",
X"F5",
X"F5",
X"EC",
X"EA",
X"E1",
X"F2",
X"FA",
X"F8",
X"0B",
X"02",
X"00",
X"FB",
X"F7",
X"D7",
X"CF",
X"CD",
X"CD",
X"CC",
X"D2",
X"D5",
X"CC",
X"E8",
X"ED",
X"F5",
X"F7",
X"FF",
X"01",
X"0A",
X"FB",
X"F2",
X"FC",
X"00",
X"1C",
X"25",
X"28",
X"2E",
X"4A",
X"4E",
X"48",
X"40",
X"38",
X"31",
X"2A",
X"1C",
X"EB",
X"DF",
X"DD",
X"D9",
X"D5",
X"D3",
X"CD",
X"DE",
X"E8",
X"DE",
X"DF",
X"D5",
X"E5",
X"F1",
X"EB",
X"D8",
X"DC",
X"E4",
X"EA",
X"F1",
X"F7",
X"FB",
X"08",
X"26",
X"18",
X"0A",
X"0F",
X"13",
X"16",
X"1D",
X"0C",
X"05",
X"0E",
X"10",
X"16",
X"10",
X"13",
X"27",
X"38",
X"32",
X"2B",
X"23",
X"1D",
X"16",
X"13",
X"00",
X"E7",
X"E8",
X"DE",
X"C4",
X"BE",
X"BD",
X"B7",
X"CC",
X"D3",
X"D1",
X"D8",
X"DE",
X"E5",
X"ED",
X"F0",
X"F4",
X"00",
X"00",
X"08",
X"0A",
X"12",
X"11",
X"25",
X"3B",
X"3A",
X"3E",
X"41",
X"30",
X"26",
X"2E",
X"10",
X"03",
X"00",
X"FC",
X"F6",
X"F3",
X"EC",
X"EE",
X"FF",
X"0A",
X"16",
X"09",
X"08",
X"00",
X"00",
X"EB",
X"D6",
X"D5",
X"D0",
X"CE",
X"D1",
X"CB",
X"BC",
X"E0",
X"EB",
X"F2",
X"F7",
X"FD",
X"00",
X"06",
X"04",
X"F4",
X"F8",
X"02",
X"20",
X"20",
X"29",
X"27",
X"3D",
X"4F",
X"4C",
X"49",
X"3F",
X"38",
X"30",
X"26",
X"EF",
X"E5",
X"E1",
X"DC",
X"D8",
X"D6",
X"D1",
X"D5",
X"EA",
X"E4",
X"E2",
X"DD",
X"F5",
X"F1",
X"F1",
X"E0",
X"D4",
X"E0",
X"E3",
X"EC",
X"F0",
X"F8",
X"FB",
X"1B",
X"0C",
X"07",
X"0F",
X"11",
X"15",
X"1B",
X"18",
X"02",
X"0C",
X"0C",
X"15",
X"10",
X"25",
X"26",
X"30",
X"3A",
X"2D",
X"2A",
X"20",
X"1C",
X"13",
X"0F",
X"EE",
X"EC",
X"D7",
X"C2",
X"C2",
X"BF",
X"BB",
X"C2",
X"D8",
X"D0",
X"D7",
X"D9",
X"E5",
X"E5",
X"FA",
X"00",
X"F6",
X"00",
X"01",
X"08",
X"0B",
X"12",
X"15",
X"35",
X"38",
X"3C",
X"39",
X"24",
X"26",
X"2C",
X"21",
X"06",
X"05",
X"FE",
X"FC",
X"F5",
X"F3",
X"EA",
X"FE",
X"1B",
X"15",
X"10",
X"09",
X"04",
X"00",
X"F9",
X"DB",
X"D6",
X"D3",
X"CF",
X"CE",
X"BC",
X"B7",
X"CE",
X"E9",
X"E8",
X"EE",
X"F3",
X"FA",
X"FE",
X"03",
X"FA",
X"F4",
X"0B",
X"19",
X"1B",
X"21",
X"22",
X"29",
X"40",
X"44",
X"41",
X"3C",
X"33",
X"2D",
X"1B",
X"FE",
X"ED",
X"EA",
X"E5",
X"E2",
X"DE",
X"DA",
X"D6",
X"E3",
X"E8",
X"DF",
X"E6",
X"F3",
X"EB",
X"E9",
X"E3",
X"D1",
X"D8",
X"E0",
X"E6",
X"EB",
X"F3",
X"F7",
X"00",
X"02",
X"03",
X"0A",
X"0E",
X"14",
X"16",
X"1C",
X"0D",
X"0C",
X"13",
X"15",
X"1B",
X"2F",
X"2B",
X"27",
X"34",
X"2B",
X"26",
X"1E",
X"1A",
X"10",
X"0E",
X"FC",
X"EA",
X"D6",
X"CC",
X"CC",
X"C6",
X"C7",
X"C1",
X"D4",
X"D5",
X"D3",
X"D6",
X"DF",
X"E2",
X"FB",
X"03",
X"F3",
X"FC",
X"FE",
X"04",
X"05",
X"0E",
X"0E",
X"22",
X"30",
X"33",
X"2A",
X"1F",
X"27",
X"27",
X"2C",
X"16",
X"0E",
X"09",
X"04",
X"FE",
X"FD",
X"F3",
X"FF",
X"1B",
X"10",
X"0D",
X"05",
X"03",
X"FC",
X"FB",
X"E7",
X"D8",
X"D6",
X"D4",
X"CA",
X"B6",
X"BE",
X"C4",
X"E1",
X"EA",
X"EF",
X"F5",
X"FC",
X"00",
X"06",
X"02",
X"FA",
X"14",
X"17",
X"1C",
X"1E",
X"24",
X"25",
X"37",
X"45",
X"43",
X"42",
X"3B",
X"34",
X"17",
X"0D",
X"F7",
X"EF",
X"EB",
X"E7",
X"E2",
X"E0",
X"DB",
X"DF",
X"EE",
X"E4",
X"F4",
X"F6",
X"F1",
X"EC",
X"EA",
X"D8",
X"D1",
X"DC",
X"E1",
X"E9",
X"ED",
X"F6",
X"ED",
X"FD",
X"04",
X"07",
X"0C",
X"10",
X"15",
X"1B",
X"17",
X"07",
X"11",
X"10",
X"23",
X"32",
X"2F",
X"28",
X"31",
X"34",
X"29",
X"24",
X"1C",
X"17",
X"0F",
X"0B",
X"EA",
X"D3",
X"D2",
X"CF",
X"CB",
X"CA",
X"C5",
X"CC",
X"DB",
X"D2",
X"D6",
X"D7",
X"E4",
X"FC",
X"02",
X"F6",
X"F4",
X"FC",
X"00",
X"04",
X"09",
X"0D",
X"14",
X"2D",
X"2F",
X"1F",
X"1F",
X"25",
X"25",
X"2D",
X"22",
X"11",
X"0F",
X"07",
X"03",
X"FF",
X"FB",
X"05",
X"19",
X"16",
X"10",
X"0A",
X"05",
X"00",
X"FC",
X"F3",
X"DB",
X"D7",
X"D5",
X"C3",
X"B5",
X"BC",
X"BD",
X"D2",
X"E6",
X"EB",
X"F2",
X"F8",
X"FE",
X"01",
X"05",
X"02",
X"10",
X"12",
X"18",
X"1B",
X"21",
X"22",
X"2C",
X"41",
X"43",
X"44",
X"41",
X"32",
X"17",
X"19",
X"08",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"01",
X"FF",
X"01",
X"FD",
X"0F",
X"2B",
X"0D",
X"09",
X"0E",
X"13",
X"1F",
X"11",
X"03",
X"16",
X"07",
X"0A",
X"14",
X"12",
X"0D",
X"0D",
X"0A",
X"0D",
X"04",
X"00",
X"0B",
X"07",
X"0D",
X"07",
X"08",
X"09",
X"04",
X"08",
X"01",
X"06",
X"0A",
X"0D",
X"10",
X"06",
X"FE",
X"FA",
X"00",
X"09",
X"09",
X"FF",
X"00",
X"08",
X"07",
X"F4",
X"07",
X"07",
X"FD",
X"FF",
X"00",
X"05",
X"08",
X"0E",
X"00",
X"01",
X"00",
X"F8",
X"FF",
X"0E",
X"02",
X"F4",
X"04",
X"FF",
X"02",
X"00",
X"F4",
X"FE",
X"FB",
X"0A",
X"FB",
X"09",
X"0C",
X"05",
X"F8",
X"06",
X"F5",
X"06",
X"06",
X"0F",
X"F3",
X"FB",
X"02",
X"FC",
X"00",
X"F5",
X"00",
X"F7",
X"00",
X"00",
X"07",
X"0B",
X"03",
X"02",
X"00",
X"F2",
X"00",
X"FD",
X"06",
X"FF",
X"08",
X"10",
X"01",
X"E5",
X"07",
X"F0",
X"00",
X"EB",
X"FC",
X"F6",
X"05",
X"F7",
X"04",
X"05",
X"00",
X"F9",
X"FC",
X"FF",
X"01",
X"03",
X"01",
X"08",
X"07",
X"FE",
X"F7",
X"00",
X"F4",
X"03",
X"FB",
X"0B",
X"FD",
X"08",
X"FD",
X"FF",
X"EA",
X"EC",
X"EA",
X"ED",
X"ED",
X"EF",
X"EF",
X"F2",
X"F0",
X"F2",
X"F1",
X"F4",
X"F3",
X"F4",
X"F3",
X"F6",
X"F5",
X"F6",
X"F6",
X"F7",
X"F7",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FD",
X"F8",
X"F4",
X"F1",
X"ED",
X"E9",
X"E6",
X"E3",
X"E0",
X"DD",
X"DA",
X"D7",
X"D5",
X"D2",
X"D0",
X"CE",
X"CB",
X"CA",
X"C7",
X"C6",
X"C9",
X"CD",
X"D5",
X"DA",
X"E1",
X"E6",
X"EC",
X"F1",
X"F6",
X"FA",
X"FF",
X"01",
X"05",
X"09",
X"0D",
X"11",
X"15",
X"18",
X"1B",
X"1E",
X"21",
X"24",
X"27",
X"2A",
X"29",
X"26",
X"1F",
X"1A",
X"14",
X"0F",
X"0A",
X"05",
X"00",
X"FE",
X"FA",
X"F6",
X"F2",
X"EF",
X"EB",
X"E8",
X"E4",
X"E1",
X"DF",
X"DC",
X"D9",
X"D6",
X"D4",
X"D1",
X"D0",
X"D4",
X"D9",
X"DF",
X"E4",
X"EA",
X"EE",
X"F4",
X"F8",
X"FD",
X"00",
X"04",
X"08",
X"0D",
X"0F",
X"13",
X"16",
X"1A",
X"1C",
X"20",
X"23",
X"27",
X"28",
X"2C",
X"2C",
X"2B",
X"25",
X"20",
X"19",
X"15",
X"0D",
X"0D",
X"02",
X"1E",
X"2D",
X"22",
X"1E",
X"18",
X"11",
X"0F",
X"FD",
X"D6",
X"D9",
X"F9",
X"00",
X"F8",
X"F8",
X"EF",
X"EE",
X"EB",
X"F1",
X"F3",
X"FD",
X"E1",
X"D3",
X"E1",
X"09",
X"13",
X"14",
X"19",
X"1C",
X"21",
X"20",
X"3A",
X"59",
X"52",
X"58",
X"55",
X"5B",
X"54",
X"5D",
X"36",
X"2C",
X"25",
X"FB",
X"FB",
X"F3",
X"F2",
X"EC",
X"E9",
X"E5",
X"E3",
X"DF",
X"DF",
X"05",
X"00",
X"11",
X"2B",
X"1D",
X"1E",
X"15",
X"12",
X"0A",
X"0D",
X"E2",
X"D1",
X"D3",
X"CF",
X"D3",
X"D6",
X"E0",
X"DD",
X"BD",
X"BE",
X"DF",
X"00",
X"FE",
X"06",
X"03",
X"0B",
X"0C",
X"13",
X"13",
X"1C",
X"0C",
X"F2",
X"F6",
X"1C",
X"2F",
X"2E",
X"33",
X"32",
X"34",
X"2C",
X"2C",
X"4F",
X"47",
X"41",
X"38",
X"32",
X"2B",
X"2A",
X"0B",
X"EA",
X"ED",
X"BF",
X"B7",
X"B7",
X"B6",
X"B6",
X"B3",
X"B3",
X"B0",
X"B2",
X"AC",
X"CB",
X"E0",
X"E4",
X"15",
X"12",
X"1C",
X"19",
X"20",
X"1F",
X"28",
X"15",
X"FB",
X"02",
X"04",
X"0B",
X"0C",
X"0F",
X"13",
X"F2",
X"E9",
X"FD",
X"20",
X"22",
X"25",
X"28",
X"29",
X"27",
X"23",
X"1D",
X"18",
X"0D",
X"ED",
X"DF",
X"F8",
X"06",
X"FF",
X"FD",
X"F6",
X"F4",
X"F1",
X"EB",
X"03",
X"0D",
X"05",
X"04",
X"FE",
X"FC",
X"F7",
X"EB",
X"C2",
X"CE",
X"B9",
X"A9",
X"B5",
X"B9",
X"C4",
X"CA",
X"D0",
X"D6",
X"DC",
X"E0",
X"F2",
X"16",
X"18",
X"40",
X"44",
X"44",
X"46",
X"48",
X"4A",
X"4C",
X"48",
X"27",
X"25",
X"27",
X"25",
X"20",
X"16",
X"17",
X"F4",
X"E2",
X"E0",
X"FC",
X"03",
X"FB",
X"FB",
X"F2",
X"F3",
X"EE",
X"EB",
X"E5",
X"E7",
X"CB",
X"B1",
X"C5",
X"DD",
X"DB",
X"D7",
X"D7",
X"D6",
X"DE",
X"DF",
X"F5",
X"17",
X"13",
X"1D",
X"1A",
X"20",
X"22",
X"24",
X"00",
X"05",
X"01",
X"E5",
X"EA",
X"F2",
X"F5",
X"FC",
X"FE",
X"03",
X"04",
X"0B",
X"0D",
X"32",
X"2F",
X"47",
X"4F",
X"42",
X"3F",
X"35",
X"2F",
X"28",
X"25",
X"02",
X"EF",
X"F2",
X"EA",
X"EA",
X"E0",
X"E5",
X"CC",
X"B2",
X"B2",
X"C1",
X"DE",
X"D2",
X"D4",
X"D0",
X"D8",
X"DC",
X"E1",
X"E4",
X"EE",
X"EC",
X"C9",
X"F0",
X"0C",
X"1F",
X"14",
X"05",
X"21",
X"16",
X"2C",
X"1D",
X"4F",
X"55",
X"4C",
X"4C",
X"55",
X"55",
X"5C",
X"43",
X"22",
X"2A",
X"14",
X"F2",
X"FC",
X"EC",
X"EA",
X"EB",
X"ED",
X"ED",
X"F2",
X"D5",
X"F5",
X"F5",
X"F3",
X"15",
X"02",
X"0D",
X"FD",
X"0B",
X"0B",
X"F7",
X"E6",
X"C6",
X"D1",
X"DF",
X"E0",
X"DE",
X"E6",
X"EB",
X"D4",
X"D1",
X"DF",
X"02",
X"04",
X"0E",
X"09",
X"1A",
X"1A",
X"20",
X"28",
X"1E",
X"17",
X"0B",
X"07",
X"25",
X"30",
X"3A",
X"30",
X"34",
X"1E",
X"1B",
X"23",
X"2C",
X"32",
X"2A",
X"21",
X"2D",
X"24",
X"11",
X"FF",
X"E2",
X"E7",
X"DB",
X"C5",
X"C8",
X"AC",
X"BB",
X"BA",
X"B1",
X"BA",
X"B1",
X"A4",
X"C0",
X"E1",
X"F1",
X"12",
X"17",
X"22",
X"17",
X"1B",
X"19",
X"23",
X"26",
X"14",
X"18",
X"01",
X"05",
X"0E",
X"0C",
X"27",
X"F4",
X"F5",
X"F3",
X"14",
X"2E",
X"29",
X"2A",
X"2A",
X"2C",
X"23",
X"0E",
X"15",
X"0A",
X"01",
X"E8",
X"0C",
X"FC",
X"ED",
X"ED",
X"E7",
X"F5",
X"DA",
X"E2",
X"DF",
X"EA",
X"DF",
X"DD",
X"DB",
X"D8",
X"D6",
X"CC",
X"B9",
X"C5",
X"C7",
X"B9",
X"BB",
X"C3",
X"C8",
X"D0",
X"D6",
X"DE",
X"E0",
X"E8",
X"EB",
X"06",
X"15",
X"2E",
X"34",
X"34",
X"38",
X"39",
X"3B",
X"3C",
X"41",
X"30",
X"1C",
X"1C",
X"15",
X"13",
X"0A",
X"09",
X"F0",
X"E1",
X"DE",
X"E7",
X"F9",
X"F1",
X"F0",
X"EC",
X"E7",
X"E5",
X"E2",
X"DF",
X"DD",
X"D7",
X"B9",
X"C4",
X"D8",
X"D1",
X"D5",
X"D9",
X"E1",
X"E4",
X"E9",
X"EE",
X"0B",
X"14",
X"14",
X"1A",
X"1C",
X"20",
X"1D",
X"09",
X"0B",
X"11",
X"02",
X"F9",
X"00",
X"02",
X"09",
X"0B",
X"10",
X"11",
X"15",
X"0C",
X"19",
X"25",
X"33",
X"36",
X"2C",
X"27",
X"20",
X"1C",
X"15",
X"12",
X"07",
X"EB",
X"EA",
X"E3",
X"E5",
X"DE",
X"DF",
X"CA",
X"B8",
X"BA",
X"B8",
X"D0",
X"D3",
X"D6",
X"DB",
X"E1",
X"E7",
X"EC",
X"F2",
X"F5",
X"FD",
X"EC",
X"EC",
X"0A",
X"09",
X"11",
X"11",
X"18",
X"18",
X"1E",
X"1C",
X"31",
X"44",
X"42",
X"45",
X"46",
X"45",
X"43",
X"26",
X"19",
X"18",
X"08",
X"F0",
X"ED",
X"E9",
X"E7",
X"E4",
X"E1",
X"DC",
X"DC",
X"D6",
X"DA",
X"EB",
X"FE",
X"04",
X"FF",
X"FC",
X"F7",
X"F4",
X"F0",
X"EC",
X"EC",
X"D8",
X"D6",
X"DE",
X"E3",
X"E9",
X"F0",
X"EC",
X"D9",
X"E4",
X"E4",
X"FF",
X"0E",
X"0E",
X"14",
X"16",
X"19",
X"1D",
X"20",
X"23",
X"28",
X"1E",
X"0D",
X"2E",
X"2E",
X"2E",
X"26",
X"21",
X"1B",
X"18",
X"0F",
X"11",
X"23",
X"1E",
X"17",
X"14",
X"0B",
X"0A",
X"F2",
X"E3",
X"E3",
X"DE",
X"C5",
X"BC",
X"BD",
X"BA",
X"BA",
X"B7",
X"B8",
X"BB",
X"C1",
X"C7",
X"E0",
X"FD",
X"11",
X"14",
X"16",
X"1A",
X"1D",
X"21",
X"22",
X"29",
X"1D",
X"0C",
X"14",
X"15",
X"1A",
X"1C",
X"1E",
X"06",
X"0B",
X"0B",
X"18",
X"2E",
X"29",
X"23",
X"1E",
X"16",
X"12",
X"0D",
X"0A",
X"03",
X"00",
X"E1",
X"F2",
X"F8",
X"F0",
X"F0",
X"EA",
X"E9",
X"E4",
X"E3",
X"DE",
X"F2",
X"F7",
X"F0",
X"F0",
X"EA",
X"F1",
X"E6",
X"DB",
X"E2",
X"E9",
X"DE",
X"D2",
X"DD",
X"DF",
X"E9",
X"EB",
X"F2",
X"F5",
X"FC",
X"FD",
X"0A",
X"26",
X"36",
X"3A",
X"3A",
X"3C",
X"3E",
X"40",
X"42",
X"3D",
X"36",
X"1A",
X"15",
X"0E",
X"0B",
X"04",
X"01",
X"EC",
X"E2",
X"E1",
X"DC",
X"ED",
X"F0",
X"E9",
X"E8",
X"E3",
X"E2",
X"DC",
X"DD",
X"D6",
X"D9",
X"C3",
X"C5",
X"D7",
X"D4",
X"DE",
X"E2",
X"EA",
X"ED",
X"F5",
X"F6",
X"04",
X"19",
X"18",
X"1E",
X"1F",
X"24",
X"20",
X"11",
X"15",
X"19",
X"17",
X"07",
X"0C",
X"0E",
X"13",
X"16",
X"17",
X"15",
X"11",
X"0A",
X"07",
X"16",
X"28",
X"25",
X"20",
X"19",
X"14",
X"0D",
X"0A",
X"03",
X"02",
X"ED",
X"E2",
X"E0",
X"DC",
X"D9",
X"D8",
X"C8",
X"BA",
X"BC",
X"B7",
X"C9",
X"DB",
X"DF",
X"E7",
X"EB",
X"F1",
X"F4",
X"FB",
X"FE",
X"03",
X"00",
X"FB",
X"11",
X"11",
X"17",
X"19",
X"1E",
X"1F",
X"23",
X"24",
X"2A",
X"3F",
X"43",
X"44",
X"42",
X"3C",
X"33",
X"18",
X"12",
X"0B",
X"08",
X"F3",
X"E8",
X"E6",
X"E3",
X"E1",
X"DE",
X"DB",
X"D7",
X"D6",
X"D2",
X"DC",
X"F7",
X"F9",
X"F5",
X"F0",
X"EE",
X"E9",
X"EA",
X"EB",
X"F2",
X"ED",
X"E2",
X"E9",
X"EE",
X"F3",
X"FA",
X"F5",
X"E8",
X"F1",
X"F3",
X"FD",
X"11",
X"17",
X"1A",
X"1D",
X"1F",
X"23",
X"25",
X"28",
X"2A",
X"2C",
X"1E",
X"2B",
X"27",
X"21",
X"1C",
X"16",
X"11",
X"0B",
X"08",
X"01",
X"0C",
X"13",
X"0A",
X"08",
X"01",
X"00",
X"E8",
X"E0",
X"DD",
X"DC",
X"CF",
X"BD",
X"BE",
X"BA",
X"BB",
X"BD",
X"C1",
X"C9",
X"D0",
X"D5",
X"DF",
X"02",
X"14",
X"17",
X"1A",
X"1C",
X"20",
X"22",
X"26",
X"29",
X"29",
X"19",
X"19",
X"1D",
X"1E",
X"24",
X"21",
X"11",
X"14",
X"14",
X"12",
X"1D",
X"22",
X"18",
X"15",
X"0D",
X"0B",
X"04",
X"02",
X"FD",
X"FD",
X"E9",
X"ED",
X"F0",
X"EA",
X"E9",
X"E4",
X"E2",
X"DE",
X"DC",
X"D8",
X"DD",
X"EB",
X"E7",
X"EC",
X"EC",
X"F6",
X"EC",
X"E5",
X"EC",
X"F2",
X"F4",
X"E5",
X"EA",
X"EF",
X"F4",
X"F9",
X"FD",
X"01",
X"04",
X"09",
X"0A",
X"27",
X"43",
X"41",
X"44",
X"44",
X"46",
X"43",
X"3F",
X"35",
X"32",
X"1C",
X"0B",
X"09",
X"02",
X"00",
X"FB",
X"E5",
X"DD",
X"DD",
X"D6",
X"DF",
X"EC",
X"D7",
X"DA",
X"DB",
X"DD",
X"DE",
X"E0",
X"E1",
X"E3",
X"E4",
X"E6",
X"E6",
X"E8",
X"E8",
X"E9",
X"EB",
X"EB",
X"EC",
X"EE",
X"EE",
X"EE",
X"EF",
X"F0",
X"F0",
X"F1",
X"F3",
X"F2",
X"F3",
X"F4",
X"F4",
X"F5",
X"F5",
X"F6",
X"F7",
X"F6",
X"F7",
X"F7",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"03",
X"12",
X"0E",
X"1C",
X"0F",
X"07",
X"19",
X"17",
X"03",
X"05",
X"15",
X"0C",
X"0A",
X"06",
X"15",
X"08",
X"0F",
X"08",
X"06",
X"1B",
X"0E",
X"FA",
X"12",
X"00",
X"0A",
X"FF",
X"0F",
X"02",
X"08",
X"0D",
X"03",
X"09",
X"0B",
X"03",
X"08",
X"07",
X"FA",
X"07",
X"08",
X"04",
X"03",
X"10",
X"0B",
X"04",
X"00",
X"FC",
X"F7",
X"0C",
X"00",
X"06",
X"FD",
X"03",
X"14",
X"0C",
X"EE",
X"FD",
X"EA",
X"00",
X"F6",
X"06",
X"F5",
X"FC",
X"03",
X"00",
X"FE",
X"FD",
X"00",
X"10",
X"08",
X"F2",
X"10",
X"06",
X"F4",
X"FA",
X"FE",
X"FB",
X"00",
X"00",
X"00",
X"02",
X"12",
X"F5",
X"02",
X"00",
X"00",
X"0A",
X"07",
X"07",
X"F2",
X"FB",
X"FC",
X"02",
X"F6",
X"00",
X"09",
X"01",
X"02",
X"FB",
X"08",
X"07",
X"0B",
X"03",
X"F8",
X"FB",
X"FD",
X"0A",
X"F4",
X"FE",
X"00",
X"FB",
X"0C",
X"F9",
X"00",
X"0A",
X"F7",
X"00",
X"FE",
X"F5",
X"02",
X"FF",
X"10",
X"03",
X"F6",
X"0C",
X"04",
X"E8",
X"0A",
X"F7",
X"F8",
X"F9",
X"FC",
X"0C",
X"F8",
X"F4",
X"07",
X"FF",
X"FD",
X"00",
X"03",
X"07",
X"03",
X"00",
X"00",
X"0A",
X"07",
X"FF",
X"00",
X"00",
X"FF",
X"04",
X"06",
X"02",
X"FC",
X"02",
X"FC",
X"00",
X"00",
X"00",
X"0A",
X"FA",
X"01",
X"FD",
X"00",
X"02",
X"F9",
X"06",
X"06",
X"04",
X"02",
X"F5",
X"FA",
X"00",
X"00",
X"01",
X"00",
X"06",
X"06",
X"FD",
X"00",
X"FD",
X"00",
X"06",
X"06",
X"F7",
X"01",
X"FE",
X"F3",
X"00",
X"FE",
X"03",
X"00",
X"0B",
X"00",
X"F7",
X"FA",
X"FD",
X"05",
X"F5",
X"0B",
X"00",
X"F1",
X"04",
X"F9",
X"02",
X"06",
X"F5",
X"00",
X"FE",
X"FC",
X"00",
X"00",
X"00",
X"FC",
X"09",
X"05",
X"02",
X"05",
X"00",
X"F6",
X"00",
X"08",
X"00",
X"F8",
X"F9",
X"01",
X"09",
X"FA",
X"FD",
X"03",
X"03",
X"FA",
X"FE",
X"0B",
X"01",
X"01",
X"F8",
X"F9",
X"08",
X"01",
X"F8",
X"01",
X"FD",
X"02",
X"07",
X"FB",
X"FD",
X"01",
X"FC",
X"F6",
X"FE",
X"05",
X"06",
X"08",
X"00",
X"05",
X"00",
X"03",
X"07",
X"0F",
X"F6",
X"FD",
X"FF",
X"F8",
X"07",
X"00",
X"02",
X"F4",
X"06",
X"FF",
X"06",
X"07",
X"03",
X"F9",
X"00",
X"FB",
X"05",
X"05",
X"04",
X"FB",
X"00",
X"F9",
X"06",
X"0E",
X"0D",
X"DF",
X"F4",
X"E2",
X"F6",
X"EB",
X"F4",
X"EC",
X"F9",
X"FD",
X"F0",
X"F7",
X"F2",
X"FF",
X"F4",
X"01",
X"F6",
X"15",
X"F7",
X"F3",
X"FA",
X"F8",
X"00",
X"F5",
X"02",
X"05",
X"09",
X"F7",
X"00",
X"05",
X"08",
X"03",
X"02",
X"15",
X"1B",
X"E9",
X"FB",
X"F7",
X"F4",
X"F5",
X"F6",
X"02",
X"EE",
X"08",
X"F4",
X"10",
X"F4",
X"02",
X"F7",
X"0A",
X"FC",
X"11",
X"01",
X"00",
X"00",
X"F9",
X"00",
X"01",
X"0A",
X"05",
X"06",
X"10",
X"07",
X"FE",
X"03",
X"00",
X"08",
X"0C",
X"17",
X"F3",
X"F3",
X"F8",
X"F2",
X"0B",
X"ED",
X"F5",
X"F3",
X"00",
X"F5",
X"FF",
X"FA",
X"0C",
X"00",
X"F8",
X"FC",
X"07",
X"06",
X"FF",
X"04",
X"0E",
X"0D",
X"FE",
X"F0",
X"FD",
X"02",
X"F7",
X"FD",
X"FE",
X"03",
X"08",
X"04",
X"FE",
X"19",
X"FD",
X"F3",
X"03",
X"F2",
X"07",
X"F7",
X"04",
X"FB",
X"FA",
X"FB",
X"07",
X"03",
X"03",
X"05",
X"09",
X"0B",
X"00",
X"08",
X"03",
X"04",
X"01",
X"0E",
X"FF",
X"00",
X"FE",
X"00",
X"F6",
X"0F",
X"00",
X"04",
X"F9",
X"07",
X"08",
X"0B",
X"FB",
X"FD",
X"ED",
X"F7",
X"F9",
X"00",
X"FC",
X"00",
X"09",
X"19",
X"E0",
X"00",
X"ED",
X"FB",
X"FA",
X"F3",
X"FF",
X"F6",
X"FE",
X"F4",
X"07",
X"F9",
X"08",
X"F4",
X"02",
X"00",
X"0B",
X"FF",
X"FC",
X"05",
X"00",
X"06",
X"00",
X"07",
X"04",
X"FC",
X"06",
X"06",
X"FC",
X"00",
X"00",
X"06",
X"08",
X"1A",
X"F9",
X"F3",
X"F5",
X"F4",
X"FB",
X"F9",
X"07",
X"EE",
X"08",
X"FA",
X"FA",
X"FA",
X"00",
X"00",
X"0B",
X"F7",
X"02",
X"0D",
X"FA",
X"01",
X"00",
X"02",
X"0A",
X"11",
X"00",
X"00",
X"F8",
X"FB",
X"07",
X"06",
X"04",
X"F5",
X"00",
X"10",
X"FC",
X"F1",
X"00",
X"F9",
X"04",
X"F4",
X"01",
X"FC",
X"0A",
X"FD",
X"05",
X"07",
X"F7",
X"00",
X"04",
X"0C",
X"02",
X"F5",
X"02",
X"00",
X"FD",
X"04",
X"FF",
X"FF",
X"03",
X"FF",
X"05",
X"0A",
X"FE",
X"05",
X"03",
X"02",
X"04",
X"0E",
X"F9",
X"F9",
X"06",
X"EF",
X"FB",
X"03",
X"FA",
X"FF",
X"F4",
X"02",
X"0B",
X"00",
X"FF",
X"09",
X"00",
X"00",
X"06",
X"00",
X"F9",
X"0B",
X"FD",
X"01",
X"0C",
X"0A",
X"EA",
X"06",
X"FA",
X"ED",
X"FC",
X"F8",
X"F4",
X"F7",
X"00",
X"02",
X"02",
X"F9",
X"08",
X"07",
X"00",
X"03",
X"FB",
X"09",
X"0E",
X"0A",
X"EE",
X"F3",
X"F3",
X"F7",
X"00",
X"F6",
X"F9",
X"FB",
X"0D",
X"F1",
X"FB",
X"F9",
X"01",
X"0B",
X"F1",
X"01",
X"02",
X"FE",
X"FD",
X"F9",
X"08",
X"0B",
X"F5",
X"02",
X"00",
X"08",
X"01",
X"F4",
X"06",
X"FC",
X"0A",
X"00",
X"05",
X"0E",
X"F4",
X"F9",
X"08",
X"F2",
X"05",
X"FA",
X"09",
X"00",
X"09",
X"FE",
X"01",
X"FF",
X"FF",
X"0E",
X"04",
X"00",
X"00",
X"FB",
X"03",
X"09",
X"12",
X"FA",
X"F7",
X"FB",
X"F5",
X"01",
X"02",
X"07",
X"F0",
X"00",
X"FB",
X"06",
X"01",
X"09",
X"0B",
X"FE",
X"E9",
X"FE",
X"FB",
X"FA",
X"F1",
X"FE",
X"FE",
X"05",
X"00",
X"F3",
X"12",
X"F8",
X"F2",
X"FF",
X"FB",
X"0C",
X"F8",
X"EF",
X"EE",
X"EB",
X"EF",
X"EE",
X"EF",
X"EF",
X"F2",
X"F0",
X"F2",
X"F2",
X"F4",
X"F3",
X"F3",
X"F4",
X"F6",
X"F5",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F9",
X"F8",
X"FA",
X"F9",
X"FA",
X"F9",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FD",
X"FE",
X"FE",
X"FF",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"06",
X"1F",
X"07",
X"1A",
X"17",
X"09",
X"0F",
X"11",
X"13",
X"13",
X"19",
X"0B",
X"0B",
X"0E",
X"07",
X"11",
X"08",
X"0C",
X"0A",
X"06",
X"16",
X"08",
X"FF",
X"10",
X"0A",
X"00",
X"04",
X"07",
X"04",
X"0D",
X"0F",
X"F0",
X"FD",
X"F5",
X"E5",
X"EB",
X"E9",
X"F8",
X"E0",
X"E8",
X"EC",
X"F2",
X"DA",
X"EE",
X"EE",
X"F5",
X"F0",
X"F9",
X"0A",
X"03",
X"08",
X"02",
X"0A",
X"1E",
X"13",
X"0E",
X"1E",
X"05",
X"1D",
X"19",
X"25",
X"21",
X"25",
X"30",
X"2B",
X"19",
X"2C",
X"2B",
X"2F",
X"39",
X"31",
X"2B",
X"2E",
X"29",
X"2A",
X"2A",
X"11",
X"17",
X"10",
X"0D",
X"17",
X"14",
X"FC",
X"F8",
X"F3",
X"F4",
X"00",
X"F5",
X"DF",
X"E7",
X"E2",
X"F6",
X"DD",
X"DB",
X"E3",
X"E7",
X"E0",
X"D4",
X"E9",
X"E9",
X"CC",
X"CD",
X"D4",
X"CD",
X"EE",
X"D7",
X"DE",
X"E5",
X"F2",
X"F0",
X"02",
X"F8",
X"FD",
X"06",
X"00",
X"0A",
X"0D",
X"03",
X"18",
X"1A",
X"24",
X"1F",
X"1D",
X"1E",
X"19",
X"22",
X"27",
X"2A",
X"2E",
X"19",
X"2C",
X"6A",
X"3C",
X"3E",
X"39",
X"33",
X"2B",
X"27",
X"22",
X"1F",
X"18",
X"15",
X"E9",
X"E2",
X"06",
X"09",
X"03",
X"00",
X"FE",
X"FA",
X"F7",
X"F5",
X"F2",
X"EE",
X"EB",
X"E9",
X"C4",
X"B5",
X"BC",
X"B4",
X"B9",
X"B2",
X"CE",
X"E7",
X"E5",
X"EB",
X"F1",
X"F2",
X"12",
X"2B",
X"28",
X"2C",
X"2B",
X"2F",
X"2D",
X"30",
X"2F",
X"35",
X"30",
X"38",
X"1F",
X"05",
X"0B",
X"E3",
X"EB",
X"EB",
X"F1",
X"F3",
X"FA",
X"FC",
X"00",
X"00",
X"13",
X"39",
X"30",
X"32",
X"29",
X"29",
X"1E",
X"1E",
X"15",
X"15",
X"0A",
X"2A",
X"2F",
X"FE",
X"00",
X"F9",
X"F9",
X"F3",
X"F4",
X"EE",
X"EE",
X"EA",
X"E9",
X"E4",
X"E8",
X"0A",
X"0C",
X"04",
X"04",
X"FE",
X"00",
X"EC",
X"C8",
X"CD",
X"D0",
X"D6",
X"DA",
X"BB",
X"B6",
X"C0",
X"C5",
X"CC",
X"CF",
X"D7",
X"DA",
X"E1",
X"E2",
X"EB",
X"EB",
X"0E",
X"24",
X"1F",
X"49",
X"54",
X"51",
X"52",
X"54",
X"51",
X"53",
X"4F",
X"56",
X"3A",
X"21",
X"27",
X"20",
X"20",
X"17",
X"17",
X"0D",
X"0E",
X"04",
X"09",
X"EA",
X"DD",
X"FD",
X"F3",
X"F3",
X"EE",
X"EE",
X"E9",
X"E9",
X"E4",
X"E6",
X"E0",
X"E2",
X"D5",
X"B2",
X"B5",
X"B2",
X"B5",
X"B2",
X"B3",
X"B4",
X"D7",
X"DE",
X"DF",
X"E4",
X"EC",
X"12",
X"16",
X"19",
X"1A",
X"1D",
X"1E",
X"23",
X"22",
X"26",
X"26",
X"29",
X"29",
X"0B",
X"04",
X"0E",
X"F8",
X"E7",
X"EF",
X"F2",
X"F6",
X"F8",
X"FE",
X"00",
X"02",
X"21",
X"34",
X"2C",
X"2F",
X"28",
X"24",
X"1E",
X"1B",
X"13",
X"12",
X"08",
X"11",
X"16",
X"FF",
X"00",
X"F9",
X"F9",
X"F5",
X"F4",
X"EF",
X"EE",
X"E9",
X"EA",
X"E1",
X"F4",
X"0A",
X"00",
X"01",
X"FC",
X"FC",
X"F5",
X"F8",
X"D4",
X"C9",
X"CC",
X"D5",
X"CE",
X"B3",
X"BF",
X"C0",
X"CA",
X"CD",
X"D7",
X"D8",
X"E1",
X"E2",
X"EA",
X"EA",
X"F7",
X"19",
X"1E",
X"1C",
X"2D",
X"4E",
X"49",
X"4B",
X"4C",
X"4B",
X"4B",
X"4D",
X"4B",
X"28",
X"25",
X"28",
X"23",
X"22",
X"1C",
X"19",
X"13",
X"11",
X"09",
X"07",
X"02",
X"FF",
X"FE",
X"FB",
X"F7",
X"F5",
X"F2",
X"EF",
X"EC",
X"EA",
X"E7",
X"DE",
X"DF",
X"C7",
X"B5",
X"B9",
X"B4",
X"B7",
X"B5",
X"B9",
X"B2",
X"C4",
X"DB",
X"DB",
X"DE",
X"F4",
X"0C",
X"09",
X"11",
X"12",
X"15",
X"14",
X"1A",
X"1A",
X"1F",
X"1E",
X"25",
X"1A",
X"01",
X"08",
X"0A",
X"0C",
X"F0",
X"F5",
X"F6",
X"FB",
X"FE",
X"02",
X"02",
X"0B",
X"2D",
X"2E",
X"30",
X"2C",
X"2D",
X"23",
X"21",
X"19",
X"18",
X"11",
X"0F",
X"04",
X"FC",
X"03",
X"FF",
X"FF",
X"F9",
X"F7",
X"F4",
X"F2",
X"EE",
X"EB",
X"EA",
X"E7",
X"FF",
X"04",
X"FE",
X"FF",
X"F8",
X"F8",
X"F0",
X"F4",
X"E5",
X"CB",
X"CC",
X"D3",
X"C1",
X"B7",
X"C3",
X"C5",
X"CE",
X"D2",
X"D9",
X"DD",
X"E3",
X"E4",
X"ED",
X"EB",
X"02",
X"1A",
X"18",
X"1D",
X"1B",
X"3A",
X"45",
X"43",
X"45",
X"46",
X"44",
X"49",
X"3C",
X"21",
X"28",
X"27",
X"27",
X"24",
X"20",
X"19",
X"18",
X"10",
X"10",
X"06",
X"0F",
X"19",
X"FC",
X"FE",
X"F8",
X"F6",
X"F2",
X"F1",
X"ED",
X"EB",
X"E8",
X"E6",
X"E2",
X"C1",
X"BE",
X"BE",
X"BE",
X"BC",
X"BC",
X"BB",
X"BB",
X"BB",
X"D5",
X"DC",
X"DB",
X"FB",
X"01",
X"04",
X"06",
X"0A",
X"0E",
X"11",
X"13",
X"15",
X"17",
X"18",
X"1E",
X"0B",
X"01",
X"0A",
X"09",
X"11",
X"02",
X"F6",
X"FD",
X"00",
X"01",
X"06",
X"06",
X"1A",
X"2D",
X"29",
X"2F",
X"29",
X"2C",
X"25",
X"22",
X"1B",
X"18",
X"10",
X"11",
X"00",
X"ED",
X"04",
X"00",
X"00",
X"FB",
X"F8",
X"F4",
X"F4",
X"EF",
X"EE",
X"E8",
X"EF",
X"02",
X"FE",
X"FC",
X"F7",
X"F6",
X"F2",
X"F1",
X"EC",
X"ED",
X"D5",
X"CD",
X"CD",
X"B9",
X"BF",
X"C4",
X"CB",
X"D0",
X"D7",
X"DB",
X"E0",
X"E5",
X"E9",
X"EC",
X"F3",
X"0C",
X"16",
X"14",
X"19",
X"18",
X"25",
X"3C",
X"3C",
X"3C",
X"3E",
X"3E",
X"42",
X"2B",
X"23",
X"27",
X"28",
X"29",
X"26",
X"24",
X"1D",
X"1B",
X"14",
X"12",
X"0A",
X"1A",
X"25",
X"04",
X"FE",
X"FB",
X"F7",
X"F4",
X"F1",
X"EE",
X"EC",
X"E9",
X"E9",
X"D9",
X"C3",
X"C8",
X"C2",
X"C3",
X"C2",
X"C3",
X"C0",
X"C2",
X"BD",
X"CA",
X"DD",
X"E5",
X"01",
X"00",
X"06",
X"08",
X"0C",
X"0F",
X"12",
X"13",
X"16",
X"18",
X"1C",
X"19",
X"02",
X"06",
X"08",
X"0A",
X"0E",
X"0F",
X"FB",
X"FC",
X"00",
X"01",
X"04",
X"09",
X"25",
X"2A",
X"2B",
X"2E",
X"2E",
X"2B",
X"29",
X"22",
X"1E",
X"18",
X"16",
X"11",
X"F9",
X"EA",
X"FD",
X"04",
X"00",
X"FE",
X"FC",
X"F8",
X"F5",
X"F1",
X"F0",
X"EB",
X"FC",
X"05",
X"FE",
X"FE",
X"F8",
X"F8",
X"F1",
X"F1",
X"EB",
X"EE",
X"E1",
X"CF",
X"C0",
X"B3",
X"BE",
X"C1",
X"CA",
X"CD",
X"D5",
X"D8",
X"E0",
X"E2",
X"E9",
X"EA",
X"F9",
X"11",
X"11",
X"16",
X"17",
X"1B",
X"1A",
X"32",
X"3D",
X"3C",
X"3E",
X"3F",
X"3B",
X"23",
X"25",
X"26",
X"29",
X"2A",
X"29",
X"26",
X"21",
X"1C",
X"18",
X"12",
X"12",
X"24",
X"25",
X"14",
X"FD",
X"FC",
X"F8",
X"F5",
X"F2",
X"EE",
X"EC",
X"E9",
X"E7",
X"CE",
X"C5",
X"C6",
X"C5",
X"C4",
X"C3",
X"C3",
X"C2",
X"C1",
X"C0",
X"C1",
X"D6",
X"F3",
X"FF",
X"00",
X"02",
X"06",
X"0A",
X"0C",
X"10",
X"12",
X"15",
X"17",
X"1B",
X"0D",
X"00",
X"07",
X"07",
X"0E",
X"0C",
X"14",
X"05",
X"FB",
X"FF",
X"00",
X"03",
X"0F",
X"23",
X"21",
X"25",
X"24",
X"2A",
X"26",
X"27",
X"21",
X"1D",
X"17",
X"14",
X"0A",
X"F5",
X"F3",
X"F2",
X"01",
X"00",
X"FD",
X"F9",
X"F6",
X"F3",
X"F1",
X"EE",
X"ED",
X"FF",
X"FD",
X"F9",
X"F6",
X"F3",
X"F1",
X"EF",
X"EC",
X"E9",
X"E6",
X"E5",
X"D4",
X"B8",
X"B9",
X"C0",
X"C6",
X"CD",
X"D2",
X"D8",
X"DC",
X"E1",
X"E7",
X"EB",
X"EE",
X"01",
X"0D",
X"0D",
X"12",
X"13",
X"18",
X"17",
X"21",
X"34",
X"36",
X"36",
X"39",
X"2B",
X"21",
X"25",
X"26",
X"28",
X"2A",
X"29",
X"28",
X"25",
X"1E",
X"1B",
X"13",
X"1A",
X"25",
X"1D",
X"1B",
X"04",
X"FB",
X"FA",
X"F6",
X"F3",
X"F0",
X"EE",
X"ED",
X"E4",
X"CE",
X"D0",
X"CC",
X"CC",
X"CA",
X"CA",
X"C7",
X"C8",
X"C5",
X"C6",
X"C1",
X"CD",
X"F4",
X"F2",
X"F9",
X"FC",
X"00",
X"01",
X"04",
X"07",
X"0A",
X"0D",
X"11",
X"13",
X"02",
X"01",
X"05",
X"08",
X"0C",
X"0E",
X"11",
X"13",
X"03",
X"02",
X"06",
X"07",
X"1C",
X"26",
X"26",
X"29",
X"29",
X"2D",
X"2C",
X"2A",
X"27",
X"21",
X"1D",
X"19",
X"06",
X"F8",
X"FA",
X"F2",
X"FE",
X"04",
X"00",
X"FE",
X"FB",
X"F8",
X"F6",
X"F0",
X"F9",
X"03",
X"FE",
X"FD",
X"F8",
X"F7",
X"F2",
X"F1",
X"EC",
X"EC",
X"E6",
X"E9",
X"D8",
X"B6",
X"B9",
X"BE",
X"C6",
X"CA",
X"D1",
X"D5",
X"DC",
X"E0",
X"E6",
X"E9",
X"F1",
X"07",
X"0B",
X"0D",
X"10",
X"13",
X"15",
X"19",
X"19",
X"2B",
X"36",
X"35",
X"38",
X"23",
X"23",
X"25",
X"27",
X"28",
X"2A",
X"2C",
X"29",
X"28",
X"22",
X"1D",
X"17",
X"25",
X"28",
X"1F",
X"1E",
X"11",
X"FE",
X"FB",
X"F8",
X"F4",
X"F2",
X"EE",
X"EE",
X"DA",
X"CF",
X"D0",
X"CD",
X"CC",
X"CB",
X"CA",
X"C9",
X"C8",
X"C7",
X"C7",
X"C4",
X"CE",
X"F0",
X"F3",
X"F6",
X"FB",
X"FD",
X"00",
X"03",
X"06",
X"09",
X"0B",
X"0F",
X"0A",
X"FD",
X"02",
X"02",
X"08",
X"09",
X"0F",
X"0E",
X"15",
X"0C",
X"00",
X"05",
X"0B",
X"23",
X"22",
X"26",
X"26",
X"29",
X"29",
X"2D",
X"29",
X"29",
X"23",
X"1F",
X"18",
X"00",
X"FC",
X"F9",
X"F6",
X"F4",
X"04",
X"FF",
X"ED",
X"EF",
X"F0",
X"F0",
X"F1",
X"F2",
X"F2",
X"F3",
X"F4",
X"F4",
X"F4",
X"F5",
X"F6",
X"F6",
X"F6",
X"F7",
X"F7",
X"F7",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"0E",
X"0C",
X"11",
X"15",
X"15",
X"0E",
X"0E",
X"10",
X"16",
X"1A",
X"0C",
X"10",
X"18",
X"06",
X"09",
X"22",
X"02",
X"F3",
X"05",
X"F6",
X"0A",
X"F6",
X"10",
X"01",
X"03",
X"FB",
X"00",
X"00",
X"09",
X"01",
X"05",
X"10",
X"0A",
X"09",
X"FD",
X"06",
X"05",
X"06",
X"0E",
X"13",
X"04",
X"04",
X"02",
X"FA",
X"04",
X"03",
X"07",
X"02",
X"05",
X"11",
X"0B",
X"F1",
X"06",
X"F3",
X"F9",
X"FA",
X"02",
X"00",
X"FC",
X"01",
X"06",
X"07",
X"EF",
X"0F",
X"F8",
X"00",
X"00",
X"05",
X"0D",
X"04",
X"F8",
X"FE",
X"F8",
X"03",
X"F8",
X"03",
X"FE",
X"09",
X"0B",
X"FD",
X"00",
X"04",
X"FE",
X"0D",
X"05",
X"EE",
X"03",
X"01",
X"00",
X"F9",
X"FA",
X"00",
X"01",
X"07",
X"00",
X"0E",
X"03",
X"F7",
X"FE",
X"03",
X"FF",
X"FE",
X"0A",
X"08",
X"F4",
X"02",
X"FF",
X"03",
X"07",
X"01",
X"FD",
X"F7",
X"04",
X"00",
X"FC",
X"FF",
X"00",
X"0B",
X"11",
X"05",
X"F0",
X"FF",
X"F4",
X"00",
X"04",
X"00",
X"F7",
X"FB",
X"08",
X"05",
X"00",
X"EC",
X"EA",
X"EB",
X"ED",
X"ED",
X"EE",
X"EE",
X"F0",
X"F0",
X"F2",
X"F1",
X"F2",
X"F2",
X"F4",
X"F4",
X"F5",
X"F4",
X"F6",
X"F5",
X"F7",
X"F7",
X"F8",
X"F7",
X"F8",
X"F8",
X"F9",
X"F9",
X"FA",
X"F9",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FD",
X"FC",
X"FD",
X"FC",
X"FD",
X"FD",
X"FE",
X"FD",
X"FE",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"07",
X"2D",
X"28",
X"2A",
X"05",
X"F7",
X"FC",
X"F9",
X"FD",
X"FA",
X"FE",
X"F9",
X"FF",
X"F7",
X"14",
X"2A",
X"24",
X"25",
X"22",
X"21",
X"21",
X"00",
X"F0",
X"F4",
X"F2",
X"F4",
X"F5",
X"F6",
X"1C",
X"20",
X"20",
X"07",
X"EC",
X"F4",
X"F0",
X"F5",
X"F4",
X"F3",
X"0F",
X"23",
X"1B",
X"20",
X"18",
X"1C",
X"15",
X"1B",
X"14",
X"1B",
X"00",
X"E7",
X"EB",
X"EF",
X"17",
X"15",
X"19",
X"FA",
X"E7",
X"EB",
X"EA",
X"EC",
X"EC",
X"ED",
X"12",
X"1B",
X"19",
X"05",
X"E5",
X"F0",
X"ED",
X"1C",
X"13",
X"1E",
X"FA",
X"EA",
X"E9",
X"F7",
X"18",
X"18",
X"16",
X"17",
X"12",
X"16",
X"00",
X"E3",
X"EA",
X"EA",
X"16",
X"14",
X"17",
X"FA",
X"E3",
X"EB",
X"E9",
X"EB",
X"ED",
X"EC",
X"0C",
X"1B",
X"14",
X"19",
X"13",
X"15",
X"10",
X"15",
X"0E",
X"17",
X"F7",
X"E3",
X"E4",
X"EE",
X"14",
X"12",
X"13",
X"10",
X"10",
X"0E",
X"0E",
X"0D",
X"0C",
X"0C",
X"0B",
X"0A",
X"0B",
X"0B",
X"09",
X"0A",
X"04",
X"DC",
X"E1",
X"DC",
X"00",
X"0D",
X"E2",
X"E4",
X"E3",
X"E5",
X"E5",
X"E7",
X"E8",
X"E9",
X"EA",
X"EC",
X"EA",
X"EC",
X"ED",
X"EF",
X"F0",
X"F0",
X"F0",
X"F2",
X"F2",
X"F3",
X"F3",
X"F3",
X"F4",
X"F5",
X"F5",
X"F6",
X"F6",
X"F7",
X"F7",
X"F7",
X"F7",
X"F7",
X"F8",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FC",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FD",
X"F8",
X"F4",
X"F0",
X"EC",
X"E9",
X"E5",
X"E2",
X"DE",
X"DB",
X"D8",
X"D5",
X"D3",
X"D0",
X"CF",
X"D2",
X"D8",
X"DF",
X"E5",
X"EA",
X"F0",
X"F5",
X"FA",
X"FF",
X"02",
X"06",
X"0A",
X"0F",
X"12",
X"16",
X"1A",
X"1D",
X"21",
X"24",
X"27",
X"29",
X"2C",
X"2D",
X"2A",
X"24",
X"1D",
X"17",
X"12",
X"0C",
X"07",
X"02",
X"FF",
X"FB",
X"F7",
X"F3",
X"EF",
X"EB",
X"E7",
X"E4",
X"E0",
X"DD",
X"DA",
X"D7",
X"D4",
X"D1",
X"D1",
X"D4",
X"DB",
X"E1",
X"E7",
X"ED",
X"F2",
X"F8",
X"FC",
X"00",
X"03",
X"08",
X"0C",
X"0F",
X"14",
X"17",
X"1B",
X"1E",
X"20",
X"25",
X"28",
X"2B",
X"2D",
X"2D",
X"2B",
X"24",
X"1D",
X"18",
X"11",
X"0E",
X"07",
X"03",
X"00",
X"FB",
X"F6",
X"F4",
X"EF",
X"EB",
X"E7",
X"E5",
X"DF",
X"1D",
X"35",
X"28",
X"27",
X"1B",
X"1A",
X"F1",
X"F3",
X"F8",
X"00",
X"00",
X"DE",
X"DD",
X"E7",
X"E7",
X"14",
X"22",
X"23",
X"26",
X"2B",
X"2B",
X"2F",
X"2F",
X"37",
X"17",
X"06",
X"2E",
X"44",
X"3C",
X"3E",
X"31",
X"30",
X"22",
X"3B",
X"4B",
X"3D",
X"39",
X"30",
X"2A",
X"24",
X"20",
X"0C",
X"CD",
X"B4",
X"B4",
X"B3",
X"B1",
X"B3",
X"AE",
X"B0",
X"AA",
X"C0",
X"E5",
X"E7",
X"EF",
X"F3",
X"FB",
X"27",
X"2B",
X"31",
X"25",
X"03",
X"0A",
X"0D",
X"13",
X"16",
X"19",
X"1D",
X"1E",
X"29",
X"53",
X"58",
X"36",
X"26",
X"2B",
X"24",
X"20",
X"19",
X"13",
X"E4",
X"DD",
X"DD",
X"DA",
X"D5",
X"D2",
X"D0",
X"CB",
X"DE",
X"1F",
X"1C",
X"1A",
X"0F",
X"0F",
X"05",
X"05",
X"FD",
X"FF",
X"D6",
X"CC",
X"D9",
X"DD",
X"E4",
X"E3",
X"BE",
X"CB",
X"C8",
X"F1",
X"09",
X"0B",
X"0D",
X"12",
X"12",
X"1C",
X"1A",
X"23",
X"0B",
X"F8",
X"FF",
X"26",
X"35",
X"33",
X"2E",
X"28",
X"1F",
X"2D",
X"46",
X"3A",
X"36",
X"2D",
X"26",
X"22",
X"18",
X"19",
X"EA",
X"AA",
X"B4",
X"AC",
X"B1",
X"AB",
X"AE",
X"AA",
X"AB",
X"AF",
X"D6",
X"D7",
X"DF",
X"E4",
X"EB",
X"F7",
X"1F",
X"1C",
X"20",
X"FE",
X"02",
X"02",
X"0C",
X"0C",
X"14",
X"13",
X"1A",
X"1C",
X"46",
X"49",
X"4D",
X"29",
X"26",
X"24",
X"24",
X"1A",
X"18",
X"F1",
X"E5",
X"E0",
X"DF",
X"DB",
X"DB",
X"D3",
X"D7",
X"CB",
X"00",
X"1E",
X"12",
X"0F",
X"07",
X"03",
X"00",
X"FB",
X"FA",
X"DE",
X"C9",
X"D1",
X"D8",
X"DE",
X"E7",
X"DF",
X"C6",
X"CE",
X"E6",
X"07",
X"04",
X"0D",
X"0C",
X"14",
X"14",
X"19",
X"1E",
X"14",
X"F8",
X"01",
X"03",
X"2F",
X"31",
X"31",
X"2B",
X"25",
X"26",
X"44",
X"37",
X"36",
X"2A",
X"27",
X"1D",
X"1D",
X"12",
X"0F",
X"C8",
X"B6",
X"B8",
X"B7",
X"B3",
X"B5",
X"B0",
X"B2",
X"B0",
X"D3",
X"D8",
X"DE",
X"E0",
X"EB",
X"EB",
X"01",
X"21",
X"21",
X"04",
X"00",
X"05",
X"0A",
X"0E",
X"12",
X"15",
X"1A",
X"1B",
X"3D",
X"4D",
X"4C",
X"49",
X"27",
X"28",
X"28",
X"21",
X"1D",
X"00",
X"E7",
X"E9",
X"E2",
X"E1",
X"DB",
X"DA",
X"D5",
X"D3",
X"DE",
X"0B",
X"0E",
X"08",
X"03",
X"00",
X"FC",
X"F9",
X"F7",
X"E4",
X"C7",
X"CF",
X"CF",
X"DA",
X"DC",
X"E9",
X"DB",
X"C9",
X"DD",
X"FE",
X"00",
X"05",
X"08",
X"0C",
X"0F",
X"15",
X"18",
X"17",
X"FE",
X"01",
X"03",
X"0E",
X"2F",
X"34",
X"30",
X"2A",
X"25",
X"3E",
X"3A",
X"33",
X"2B",
X"26",
X"1E",
X"1A",
X"13",
X"0E",
X"EE",
X"C8",
X"BD",
X"BE",
X"BA",
X"BC",
X"B8",
X"B8",
X"B3",
X"CD",
X"D8",
X"D6",
X"DC",
X"E2",
X"EA",
X"EC",
X"01",
X"1F",
X"05",
X"FE",
X"01",
X"07",
X"0A",
X"10",
X"11",
X"17",
X"15",
X"2E",
X"46",
X"41",
X"48",
X"3E",
X"25",
X"2A",
X"25",
X"25",
X"0E",
X"F2",
X"F2",
X"ED",
X"E9",
X"E7",
X"E2",
X"E1",
X"D9",
X"E2",
X"FB",
X"0F",
X"12",
X"09",
X"06",
X"00",
X"FD",
X"FB",
X"F0",
X"CE",
X"CD",
X"CF",
X"D5",
X"DB",
X"E1",
X"EB",
X"D9",
X"CF",
X"FB",
X"FD",
X"04",
X"04",
X"0C",
X"0D",
X"13",
X"15",
X"1A",
X"00",
X"00",
X"04",
X"08",
X"14",
X"37",
X"31",
X"34",
X"28",
X"42",
X"3C",
X"2C",
X"26",
X"22",
X"19",
X"16",
X"0D",
X"0D",
X"F3",
X"E3",
X"C8",
X"C3",
X"C1",
X"C0",
X"BC",
X"BD",
X"B7",
X"C9",
X"D4",
X"D1",
X"D4",
X"DA",
X"E0",
X"E8",
X"E9",
X"05",
X"07",
X"F6",
X"00",
X"01",
X"07",
X"0A",
X"0E",
X"13",
X"14",
X"23",
X"3C",
X"3A",
X"3E",
X"40",
X"36",
X"23",
X"2A",
X"26",
X"1B",
X"FC",
X"FD",
X"F4",
X"F4",
X"ED",
X"EC",
X"E6",
X"E4",
X"E2",
X"FA",
X"F7",
X"0D",
X"06",
X"03",
X"FE",
X"FD",
X"F6",
X"F3",
X"D3",
X"D0",
X"CC",
X"D2",
X"D5",
X"E0",
X"E0",
X"EC",
X"D7",
X"EE",
X"FB",
X"FF",
X"00",
X"07",
X"08",
X"10",
X"10",
X"19",
X"04",
X"00",
X"05",
X"0C",
X"0B",
X"20",
X"34",
X"33",
X"2D",
X"3A",
X"42",
X"36",
X"31",
X"29",
X"23",
X"1E",
X"16",
X"15",
X"00",
X"EB",
X"E7",
X"C9",
X"C9",
X"C5",
X"C4",
X"C0",
X"BD",
X"C6",
X"DB",
X"D2",
X"D5",
X"D5",
X"DD",
X"E1",
X"E9",
X"EE",
X"03",
X"F6",
X"FE",
X"00",
X"05",
X"08",
X"0D",
X"10",
X"15",
X"1C",
X"3A",
X"39",
X"3F",
X"3D",
X"44",
X"32",
X"27",
X"2A",
X"24",
X"04",
X"00",
X"FB",
X"F8",
X"F2",
X"F0",
X"EA",
X"E8",
X"E2",
X"FA",
X"F8",
X"FB",
X"0C",
X"05",
X"01",
X"FF",
X"F9",
X"F8",
X"DC",
X"D0",
X"D1",
X"D0",
X"D3",
X"DA",
X"DF",
X"E7",
X"E8",
X"EA",
X"F7",
X"FA",
X"FF",
X"02",
X"07",
X"0B",
X"0E",
X"15",
X"08",
X"FD",
X"05",
X"05",
X"0C",
X"0C",
X"24",
X"36",
X"2E",
X"3B",
X"46",
X"3C",
X"37",
X"2F",
X"29",
X"22",
X"1C",
X"18",
X"0A",
X"EF",
X"F1",
X"E0",
X"C9",
X"C8",
X"C5",
X"C4",
X"C0",
X"C5",
X"DA",
X"D6",
X"D5",
X"D3",
X"D7",
X"DE",
X"E3",
X"E9",
X"EE",
X"F3",
X"FA",
X"FD",
X"01",
X"05",
X"09",
X"0C",
X"12",
X"14",
X"31",
X"39",
X"3A",
X"3D",
X"3E",
X"41",
X"30",
X"25",
X"2B",
X"0E",
X"02",
X"00",
X"FC",
X"F6",
X"F4",
X"EE",
X"EC",
X"E5",
X"F6",
X"00",
X"F5",
X"FF",
X"0C",
X"02",
X"01",
X"FB",
X"FB",
X"E4",
X"D2",
X"D2",
X"CE",
X"CF",
X"D4",
X"D8",
X"E1",
X"E4",
X"F5",
X"F4",
X"F6",
X"FD",
X"00",
X"03",
X"08",
X"0B",
X"11",
X"0A",
X"FB",
X"00",
X"03",
X"07",
X"0E",
X"0F",
X"25",
X"2F",
X"31",
X"41",
X"37",
X"32",
X"2A",
X"25",
X"1E",
X"18",
X"13",
X"0A",
X"F3",
X"EE",
X"ED",
X"DE",
X"CB",
X"CD",
X"C7",
X"C8",
X"C4",
X"D9",
X"D7",
X"D4",
X"D1",
X"D3",
X"D5",
X"DE",
X"E2",
X"E9",
X"DE",
X"F3",
X"F8",
X"FF",
X"00",
X"06",
X"07",
X"0E",
X"0F",
X"25",
X"30",
X"32",
X"33",
X"38",
X"37",
X"3C",
X"29",
X"29",
X"1A",
X"0B",
X"07",
X"03",
X"00",
X"FD",
X"F6",
X"F4",
X"ED",
X"F6",
X"00",
X"FB",
X"F5",
X"FE",
X"04",
X"FF",
X"FC",
X"F6",
X"EB",
X"D5",
X"D5",
X"D1",
X"CF",
X"D1",
X"D5",
X"DB",
X"E1",
X"EE",
X"00",
X"EF",
X"F8",
X"FB",
X"00",
X"02",
X"09",
X"0C",
X"0D",
X"FD",
X"02",
X"04",
X"0C",
X"0D",
X"14",
X"15",
X"2E",
X"34",
X"48",
X"43",
X"3C",
X"33",
X"2E",
X"25",
X"22",
X"1A",
X"15",
X"FC",
X"F6",
X"F0",
X"F0",
X"DB",
X"CF",
X"CD",
X"CB",
X"C7",
X"D7",
X"DC",
X"D8",
X"D5",
X"D3",
X"D3",
X"DA",
X"DE",
X"E8",
X"DA",
X"DF",
X"F9",
X"FB",
X"00",
X"03",
X"08",
X"0B",
X"0E",
X"1F",
X"2F",
X"2F",
X"33",
X"34",
X"37",
X"39",
X"3A",
X"29",
X"1F",
X"0F",
X"0E",
X"06",
X"04",
X"00",
X"FC",
X"F6",
X"F1",
X"F6",
X"02",
X"FC",
X"FB",
X"F3",
X"00",
X"02",
X"FE",
X"FB",
X"F1",
X"DA",
X"D8",
X"D3",
X"D3",
X"D0",
X"D2",
X"D5",
X"DD",
X"E4",
X"00",
X"FB",
X"F2",
X"F8",
X"FC",
X"00",
X"04",
X"08",
X"0C",
X"FD",
X"FF",
X"02",
X"07",
X"0B",
X"10",
X"13",
X"1A",
X"30",
X"45",
X"49",
X"41",
X"39",
X"32",
X"2C",
X"25",
X"1F",
X"1A",
X"04",
X"F7",
X"F6",
X"F0",
X"EE",
X"D8",
X"CE",
X"CF",
X"C9",
X"D6",
X"DF",
X"D9",
X"D8",
X"D3",
X"D2",
X"D4",
X"D9",
X"E1",
X"DC",
X"D1",
X"E6",
X"F8",
X"FC",
X"00",
X"02",
X"08",
X"0A",
X"18",
X"2C",
X"2D",
X"31",
X"32",
X"35",
X"37",
X"3A",
X"38",
X"21",
X"12",
X"11",
X"0C",
X"07",
X"03",
X"FF",
X"FB",
X"F6",
X"F5",
X"03",
X"00",
X"FD",
X"F9",
X"F4",
X"01",
X"01",
X"FD",
X"F8",
X"E0",
X"DA",
X"D7",
X"D5",
X"D2",
X"D0",
X"D2",
X"D8",
X"DF",
X"F6",
X"02",
X"F7",
X"F2",
X"F2",
X"DD",
X"DF",
X"DF",
X"E1",
X"E2",
X"E4",
X"E5",
X"E6",
X"E7",
X"E8",
X"E9",
X"EA",
X"EB",
X"EC",
X"ED",
X"EE",
X"EF",
X"EF",
X"F0",
X"F1",
X"F1",
X"F2",
X"F3",
X"F3",
X"F4",
X"F4",
X"F5",
X"F5",
X"F6",
X"F6",
X"F7",
X"F7",
X"F8",
X"F8",
X"F8",
X"F9",
X"F9",
X"F9",
X"FA",
X"FA",
X"FA",
X"FA",
X"FB",
X"FB",
X"FB",
X"FB",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FC",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"01",
X"FE",
X"00",
X"FE",
X"01",
X"FF",
X"19",
X"16",
X"15",
X"15",
X"18",
X"1F",
X"1B",
X"00",
X"08",
X"05",
X"0D",
X"15",
X"F9",
X"0A",
X"00",
X"0D",
X"03",
X"15",
X"0C",
X"08",
X"07",
X"07",
X"04",
X"05",
X"03",
X"0E",
X"0D",
X"11",
X"08",
X"06",
X"00",
X"0A",
X"0B",
X"1A",
X"F3",
X"00",
X"00",
X"F9",
X"FC",
X"00",
X"12",
X"EF",
X"01",
X"F9",
X"03",
X"00",
X"00",
X"04",
X"05",
X"00",
X"05",
X"0D",
X"07",
X"03",
X"FF",
X"05",
X"0B",
X"10",
X"03",
X"F4",
X"F8",
X"F3",
X"05",
X"F9",
X"03",
X"FC",
X"08",
X"0E",
X"F2",
X"FD",
X"FC",
X"FE",
X"08",
X"01",
X"00",
X"FD",
X"FD",
X"FD",
X"FE",
X"06",
X"05",
X"0E",
X"0B",
X"00",
X"F8",
X"F9",
X"00",
X"FF",
X"08",
X"FB",
X"00",
X"08",
X"09",
X"F3",
X"10",
X"FF",
X"F1",
X"FD",
X"F7",
X"00",
X"FD",
X"0B",
X"03",
X"FB",
X"03",
X"F5",
X"FF",
X"01",
X"00",
X"02",
X"03",
X"06",
X"10",
X"FA",
X"F3",
X"00",
X"FA",
X"03",
X"EE",
X"07",
X"F7",
X"00",
X"FC",
X"04",
X"07",
X"0E",
X"FE",
X"F5",
X"07",
X"EF",
X"E8",
X"EE",
X"EC",
X"EF",
X"EF",
X"F0",
X"EF",
X"F2",
X"F2",
X"F1",
X"F3",
X"F4",
X"F3",
X"F5",
X"F5",
X"F4",
X"F6",
X"F5",
X"F6",
X"F8",
X"F7",
X"F8",
X"F8",
X"FA",
X"F8",
X"F8",
X"F9",
X"FA",
X"FA",
X"FA",
X"FB",
X"FA",
X"FB",
X"FB",
X"FC",
X"FB",
X"FD",
X"FC",
X"FD",
X"FD",
X"FC",
X"FD",
X"FD",
X"FE",
X"FD",
X"FD",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FE",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"FF",
X"FF",
X"FF",
X"00",
X"00",
X"00",
X"FF",
X"00",
X"FF",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"06",
X"0B",
X"0F",
X"14",
X"18",
X"1C",
X"20",
X"24",
X"27",
X"2A",
X"2E",
X"31",
X"34",
X"35",
X"32",
X"2B",
X"24",
X"1D",
X"17",
X"11",
X"0B",
X"05",
X"00",
X"FD",
X"F8",
X"F3",
X"EE",
X"EA",
X"E6",
X"E2",
X"DE",
X"DA",
X"D7",
X"D4",
X"D4",
X"D9",
X"E1",
X"E7",
X"ED",
X"F3",
X"F9",
X"FE",
X"01",
X"07",
X"0B",
X"10",
X"14",
X"19",
X"1D",
X"21",
X"24",
X"28",
X"2B",
X"2F",
X"30",
X"30",
X"30"
	);
--//--------------------------------------
  begin

    if (RESET_N='0') then
      Q <= sqr_table(0);
    elsif(rising_edge(CLK)) then
      if (ENA='1') then
          Q <= sqr_table(to_integer(unsigned(ADDR)));
      end if;
    end if;
  end process;
end arch;